CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 760 30 100 10
176 80 1918 1019
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
0 4 0.500000 0.500000
344 176 457 273
42991634 0
0
6 Title:
5 Name:
0
0
0
97
13 Logic Switch~
5 322 921 0 1 11
0 7
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V3
-7 -26 7 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
6616 0 0
2
44287.7 0
0
13 Logic Switch~
5 805 214 0 10 11
0 83 0 0 0 0 0 0 0 0
1
0
0 0 21360 270
2 5V
-6 -21 8 -13
7 VSinal2
-23 -31 26 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
365 0 0
2
44287.7 1
0
13 Logic Switch~
5 530 217 0 10 11
0 84 0 0 0 0 0 0 0 0
1
0
0 0 21360 270
2 5V
-6 -21 8 -13
7 VSinal1
-23 -31 26 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
8135 0 0
2
44287.7 1
0
13 Logic Switch~
5 950 221 0 10 11
0 85 0 0 0 0 0 0 0 0
1
0
0 0 21360 270
2 5V
-6 -21 8 -13
2 V8
-6 -31 8 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -2 0
1 V
9162 0 0
2
44287.7 6
0
13 Logic Switch~
5 917 221 0 10 11
0 86 0 0 0 0 0 0 0 0
1
0
0 0 21360 270
2 5V
-6 -21 8 -13
2 V9
-6 -31 8 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -2 0
1 V
8373 0 0
2
44287.7 4
0
13 Logic Switch~
5 883 219 0 1 11
0 87
0
0 0 21360 270
2 0V
-6 -21 8 -13
3 V10
-9 -31 12 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
5507 0 0
2
44287.7 2
0
13 Logic Switch~
5 848 218 0 1 11
0 88
0
0 0 21360 270
2 0V
-6 -21 8 -13
3 V11
-9 -31 12 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
3304 0 0
2
44287.7 0
0
13 Logic Switch~
5 302 293 0 10 11
0 80 0 0 0 0 0 0 0 0
1
0
0 0 21360 692
2 5V
-7 -16 7 -8
2 V7
-7 -26 7 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -2 0
1 V
5515 0 0
2
44287.7 0
0
13 Logic Switch~
5 680 220 0 10 11
0 97 0 0 0 0 0 0 0 0
1
0
0 0 21360 270
2 5V
-6 -21 8 -13
2 V6
-6 -31 8 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
3399 0 0
2
44287.7 0
0
13 Logic Switch~
5 647 220 0 10 11
0 98 0 0 0 0 0 0 0 0
1
0
0 0 21360 270
2 5V
-6 -21 8 -13
2 V5
-6 -31 8 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
3772 0 0
2
44287.7 0
0
13 Logic Switch~
5 613 218 0 10 11
0 99 0 0 0 0 0 0 0 0
1
0
0 0 21360 270
2 5V
-6 -21 8 -13
2 V4
-6 -31 8 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -2 0
1 V
3517 0 0
2
44287.7 0
0
13 Logic Switch~
5 578 217 0 1 11
0 100
0
0 0 21360 270
2 0V
-6 -21 8 -13
2 V1
-6 -31 8 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -2 0
1 V
6794 0 0
2
44287.7 0
0
13 Quad 3-State~
48 1031 590 0 9 19
0 65 64 63 62 39 38 37 36 52
0
0 0 4720 270
8 QUAD3STA
-28 -44 28 -36
3 U12
42 -1 63 7
0
15 DVCC=16;DGND=8;
85 %D [%16bi %8bi %1i %2i %3i %4i %9i]
+ [%16bo %1o %2o %3o %4o %9o %5o %6o %7o %8o] %M
0
12 type:digital
5 DIP16
19

0 1 2 3 4 5 6 7 8 9
1 2 3 4 5 6 7 8 9 0
65 0 0 0 1 0 0 0
1 U
7741 0 0
2
44287.7 0
0
13 Quad 3-State~
48 649 587 0 9 19
0 73 72 71 70 47 46 45 44 53
0
0 0 4720 270
8 QUAD3STA
-28 -44 28 -36
2 U7
45 -1 59 7
0
15 DVCC=16;DGND=8;
85 %D [%16bi %8bi %1i %2i %3i %4i %9i]
+ [%16bo %1o %2o %3o %4o %9o %5o %6o %7o %8o] %M
0
12 type:digital
5 DIP16
19

0 1 2 3 4 5 6 7 8 9
1 2 3 4 5 6 7 8 9 0
65 0 0 0 1 0 0 0
1 U
9229 0 0
2
44287.7 0
0
12 Quad D Flop~
47 886 404 0 9 19
0 92 91 90 89 65 64 63 62 82
0
0 0 4720 270
4 QDFF
-14 -44 14 -36
2 U5
40 -4 54 4
0
15 DVCC=16;DGND=8;
85 %D [%16bi %8bi %1i %2i %3i %4i %9i]
+ [%16bo %1o %2o %3o %4o %9o %5o %6o %7o %8o] %M
0
11 typeDigital
5 DIP16
19

0 1 2 3 4 5 6 7 8 9
1 2 3 4 5 6 7 8 9 0
65 0 0 0 1 0 0 0
1 U
5474 0 0
2
44287.7 0
0
12 Quad D Flop~
47 627 409 0 9 19
0 96 95 94 93 73 72 71 70 82
0
0 0 4720 270
4 QDFF
-14 -44 14 -36
2 U4
40 -4 54 4
0
15 DVCC=16;DGND=8;
85 %D [%16bi %8bi %1i %2i %3i %4i %9i]
+ [%16bo %1o %2o %3o %4o %9o %5o %6o %7o %8o] %M
0
11 typeDigital
5 DIP16
19

0 1 2 3 4 5 6 7 8 9
1 2 3 4 5 6 7 8 9 0
65 0 0 0 1 0 0 0
1 U
6991 0 0
2
44287.7 0
0
13 Quad 3-State~
48 883 301 0 9 19
0 85 86 87 88 92 91 90 89 81
0
0 0 4720 270
8 QUAD3STA
-28 -44 28 -36
2 U6
45 -1 59 7
0
15 DVCC=16;DGND=8;
85 %D [%16bi %8bi %1i %2i %3i %4i %9i]
+ [%16bo %1o %2o %3o %4o %9o %5o %6o %7o %8o] %M
0
12 type:digital
5 DIP16
19

0 1 2 3 4 5 6 7 8 9
1 2 3 4 5 6 7 8 9 0
65 0 0 0 1 0 0 0
1 U
4824 0 0
2
44287.7 0
0
13 Quad 3-State~
48 624 305 0 9 19
0 97 98 99 100 96 95 94 93 81
0
0 0 4720 270
8 QUAD3STA
-28 -44 28 -36
3 U11
42 -1 63 7
0
15 DVCC=16;DGND=8;
85 %D [%16bi %8bi %1i %2i %3i %4i %9i]
+ [%16bo %1o %2o %3o %4o %9o %5o %6o %7o %8o] %M
0
12 type:digital
5 DIP16
19

0 1 2 3 4 5 6 7 8 9
1 2 3 4 5 6 7 8 9 0
65 0 0 0 1 0 0 0
1 U
3594 0 0
2
44287.7 0
0
14 Logic Display~
6 363 1430 0 1 2
10 2
0
0 0 53856 180
6 100MEG
3 -16 45 -8
3 L28
11 0 32 8
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
3206 0 0
2
44287.7 0
0
5 4030~
219 360 1387 0 3 22
0 4 3 2
0
0 0 624 270
4 4030
-7 -24 21 -16
4 U23A
-12 -4 16 4
0
15 DVDD=14;DGND=7;
49 %D [%14bi %7bi %1i %2i]
+ [%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 1 15 0
1 U
9162 0 0
2
44287.7 0
0
14 Logic Display~
6 1232 1102 0 1 2
10 5
0
0 0 53856 270
6 100MEG
3 -16 45 -8
3 L27
-9 -15 12 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
9381 0 0
2
44287.7 0
0
14 Logic Display~
6 1161 1100 0 1 2
10 6
0
0 0 53856 90
6 100MEG
3 -16 45 -8
3 L26
-13 -15 8 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
4992 0 0
2
44287.7 0
0
14 Logic Display~
6 1237 1416 0 1 2
10 9
0
0 0 53856 180
6 100MEG
3 -16 45 -8
3 L25
11 0 32 8
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
8456 0 0
2
44287.7 0
0
14 Logic Display~
6 1021 1100 0 1 2
10 10
0
0 0 53856 270
6 100MEG
3 -16 45 -8
3 L24
-9 -15 12 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
8342 0 0
2
44287.7 0
0
14 Logic Display~
6 971 1102 0 1 2
10 11
0
0 0 53856 90
6 100MEG
3 -16 45 -8
3 L23
-13 -15 8 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
9685 0 0
2
44287.7 0
0
14 Logic Display~
6 1036 1184 0 1 2
10 12
0
0 0 53856 0
6 100MEG
3 -16 45 -8
3 L22
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
7318 0 0
2
44287.7 0
0
14 Logic Display~
6 1047 1411 0 1 2
10 13
0
0 0 53856 180
6 100MEG
3 -16 45 -8
3 L21
11 0 32 8
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
3167 0 0
2
44287.7 0
0
14 Logic Display~
6 841 1178 0 1 2
10 15
0
0 0 53856 0
6 100MEG
3 -16 45 -8
3 L20
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
3547 0 0
2
44287.7 0
0
14 Logic Display~
6 832 1414 0 1 2
10 18
0
0 0 53856 180
6 100MEG
3 -16 45 -8
3 L19
11 0 32 8
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
9895 0 0
2
44287.7 0
0
14 Logic Display~
6 807 1102 0 1 2
10 16
0
0 0 53856 270
6 100MEG
3 -16 45 -8
3 L18
-9 -15 12 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
5891 0 0
2
44287.7 0
0
14 Logic Display~
6 753 1103 0 1 2
10 17
0
0 0 53856 90
6 100MEG
3 -16 45 -8
3 L17
-13 -15 8 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
8863 0 0
2
44287.7 0
0
14 Logic Display~
6 610 1100 0 1 2
10 21
0
0 0 53856 270
6 100MEG
3 -16 45 -8
3 L16
-9 -15 12 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
393 0 0
2
44287.7 0
0
14 Logic Display~
6 522 1103 0 1 2
10 22
0
0 0 53856 90
6 100MEG
3 -16 45 -8
3 L15
-13 -15 8 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
6476 0 0
2
44287.7 0
0
14 Logic Display~
6 601 1414 0 1 2
10 20
0
0 0 53856 180
6 100MEG
3 -16 45 -8
3 L14
11 0 32 8
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
4421 0 0
2
44287.7 0
0
14 Logic Display~
6 621 1176 0 1 2
10 4
0
0 0 53856 0
6 100MEG
3 -16 45 -8
3 L13
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
5341 0 0
2
44287.7 0
0
5 4030~
219 1234 1373 0 3 22
0 7 8 9
0
0 0 624 270
4 4030
-7 -24 21 -16
4 U21D
-16 -7 12 1
0
15 DVDD=14;DGND=7;
49 %D [%14bi %7bi %1i %2i]
+ [%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 4 13 0
1 U
6395 0 0
2
44287.7 4
0
5 4030~
219 1182 1281 0 3 22
0 5 6 8
0
0 0 624 270
4 4030
-7 -24 21 -16
4 U21C
-12 -4 16 4
0
15 DVDD=14;DGND=7;
49 %D [%14bi %7bi %1i %2i]
+ [%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 8 9 10 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 3 13 0
1 U
8741 0 0
2
44287.7 3
0
5 4071~
219 1067 1201 0 3 22
0 25 24 12
0
0 0 624 512
4 4071
-7 -24 21 -16
4 U22A
-17 -6 11 2
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 1 14 0
1 U
8261 0 0
2
44287.7 2
0
5 4081~
219 1134 1182 0 3 22
0 6 5 25
0
0 0 624 512
4 4081
-7 -24 21 -16
4 U20D
-12 -11 16 -3
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 4 12 0
1 U
7839 0 0
2
44287.7 1
0
5 4081~
219 1135 1226 0 3 22
0 7 8 24
0
0 0 624 512
4 4081
-7 -24 21 -16
4 U20C
-13 -12 15 -4
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 8 9 10 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 3 12 0
1 U
8885 0 0
2
44287.7 0
0
5 4030~
219 1044 1368 0 3 22
0 12 14 13
0
0 0 624 270
4 4030
-7 -24 21 -16
4 U21B
-16 -7 12 1
0
15 DVDD=14;DGND=7;
49 %D [%14bi %7bi %1i %2i]
+ [%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 5 6 4 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 2 13 0
1 U
3689 0 0
2
44287.7 4
0
5 4030~
219 992 1276 0 3 22
0 10 11 14
0
0 0 624 270
4 4030
-7 -24 21 -16
4 U21A
-12 -4 16 4
0
15 DVDD=14;DGND=7;
49 %D [%14bi %7bi %1i %2i]
+ [%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 1 13 0
1 U
3570 0 0
2
44287.7 3
0
5 4071~
219 877 1196 0 3 22
0 27 26 15
0
0 0 624 512
4 4071
-7 -24 21 -16
4 U18D
-17 -6 11 2
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 4 8 0
1 U
9343 0 0
2
44287.7 2
0
5 4081~
219 931 1177 0 3 22
0 11 10 27
0
0 0 624 512
4 4081
-7 -24 21 -16
4 U20B
-12 -11 16 -3
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 5 6 4 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 2 12 0
1 U
9817 0 0
2
44287.7 1
0
5 4081~
219 933 1221 0 3 22
0 12 14 26
0
0 0 624 512
4 4081
-7 -24 21 -16
4 U20A
-13 -12 15 -4
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 1 12 0
1 U
9129 0 0
2
44287.7 0
0
5 4081~
219 714 1220 0 3 22
0 15 19 28
0
0 0 624 512
4 4081
-7 -24 21 -16
3 U1C
-10 -12 11 -4
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 8 9 10 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 3 9 0
1 U
5573 0 0
2
44287.7 2
0
5 4081~
219 716 1175 0 3 22
0 17 16 29
0
0 0 624 512
4 4081
-7 -24 21 -16
3 U1D
-9 -11 12 -3
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 4 9 0
1 U
8151 0 0
2
44287.7 1
0
5 4071~
219 659 1194 0 3 22
0 29 28 4
0
0 0 624 512
4 4071
-7 -24 21 -16
4 U18C
-17 -6 11 2
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 8 9 10 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 3 8 0
1 U
6375 0 0
2
44287.7 0
0
5 4030~
219 777 1274 0 3 22
0 16 17 19
0
0 0 624 270
4 4030
-7 -24 21 -16
4 U19D
-12 -4 16 4
0
15 DVDD=14;DGND=7;
49 %D [%14bi %7bi %1i %2i]
+ [%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 4 11 0
1 U
3122 0 0
2
44287.7 1
0
5 4030~
219 829 1366 0 3 22
0 15 19 18
0
0 0 624 270
4 4030
-7 -24 21 -16
4 U19C
-16 -7 12 1
0
15 DVDD=14;DGND=7;
49 %D [%14bi %7bi %1i %2i]
+ [%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 8 9 10 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 3 11 0
1 U
5719 0 0
2
44287.7 0
0
5 4071~
219 428 1190 0 3 22
0 31 30 3
0
0 0 624 512
4 4071
-7 -24 21 -16
4 U18B
-17 -6 11 2
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 5 6 4 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 2 8 0
1 U
3569 0 0
2
44287.7 5
0
5 4081~
219 495 1171 0 3 22
0 22 21 31
0
0 0 624 512
4 4081
-7 -24 21 -16
3 U1A
-9 -11 12 -3
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 1 9 0
1 U
7688 0 0
2
44287.7 4
0
5 4081~
219 496 1215 0 3 22
0 4 23 30
0
0 0 624 512
4 4081
-7 -24 21 -16
3 U1B
-10 -12 11 -4
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 5 6 4 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 2 9 0
1 U
3316 0 0
2
44287.7 3
0
14 Logic Display~
6 376 1163 0 1 2
10 3
0
0 0 53856 0
6 100MEG
3 -16 45 -8
3 L12
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
6741 0 0
2
44287.7 2
0
5 4030~
219 544 1278 0 3 22
0 21 22 23
0
0 0 624 270
4 4030
-7 -24 21 -16
4 U19A
-12 -4 16 4
0
15 DVDD=14;DGND=7;
49 %D [%14bi %7bi %1i %2i]
+ [%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 1 11 0
1 U
593 0 0
2
44287.7 1
0
5 4030~
219 598 1366 0 3 22
0 4 23 20
0
0 0 624 270
4 4030
-7 -24 21 -16
4 U19B
-12 -4 16 4
0
15 DVDD=14;DGND=7;
49 %D [%14bi %7bi %1i %2i]
+ [%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 5 6 4 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 2 11 0
1 U
4132 0 0
2
44287.7 0
0
5 4030~
219 1213 1029 0 3 22
0 7 35 5
0
0 0 624 270
4 4030
-7 -24 21 -16
3 U2D
-9 -4 12 4
0
15 DVDD=14;DGND=7;
49 %D [%14bi %7bi %1i %2i]
+ [%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 4 10 0
1 U
3574 0 0
2
44287.7 0
0
5 4030~
219 988 1029 0 3 22
0 7 34 10
0
0 0 624 270
4 4030
-7 -24 21 -16
3 U2C
-9 -4 12 4
0
15 DVDD=14;DGND=7;
49 %D [%14bi %7bi %1i %2i]
+ [%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 8 9 10 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 3 10 0
1 U
315 0 0
2
44287.7 0
0
5 4030~
219 796 1030 0 3 22
0 7 33 16
0
0 0 624 270
4 4030
-7 -24 21 -16
3 U2B
-9 -4 12 4
0
15 DVDD=14;DGND=7;
49 %D [%14bi %7bi %1i %2i]
+ [%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 5 6 4 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 2 10 0
1 U
3889 0 0
2
44287.7 0
0
5 4030~
219 591 1028 0 3 22
0 7 32 21
0
0 0 624 270
4 4030
-7 -24 21 -16
3 U2A
-9 -4 12 4
0
15 DVDD=14;DGND=7;
49 %D [%14bi %7bi %1i %2i]
+ [%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 1 10 0
1 U
3545 0 0
2
44287.7 2
0
5 4071~
219 1032 829 0 3 22
0 39 40 35
0
0 0 624 270
4 4071
-7 -24 21 -16
4 U18A
-9 -6 19 2
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 1 8 0
1 U
8315 0 0
2
44287.7 3
0
5 4071~
219 998 829 0 3 22
0 38 41 34
0
0 0 624 270
4 4071
-7 -24 21 -16
4 U16D
-9 -6 19 2
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 4 7 0
1 U
817 0 0
2
44287.7 2
0
5 4071~
219 965 829 0 3 22
0 37 42 33
0
0 0 624 270
4 4071
-7 -24 21 -16
4 U16C
-9 -6 19 2
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 8 9 10 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 3 7 0
1 U
9586 0 0
2
44287.7 1
0
5 4071~
219 931 829 0 3 22
0 36 43 32
0
0 0 624 270
4 4071
-7 -24 21 -16
4 U16B
-9 -6 19 2
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 5 6 4 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 2 7 0
1 U
3736 0 0
2
44287.7 0
0
5 4071~
219 651 809 0 3 22
0 47 48 6
0
0 0 624 270
4 4071
-7 -24 21 -16
4 U16A
-9 -6 19 2
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 1 7 0
1 U
4344 0 0
2
44287.7 3
0
5 4071~
219 617 809 0 3 22
0 46 49 11
0
0 0 624 270
4 4071
-7 -24 21 -16
3 U3D
-6 -6 15 2
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 4 3 0
1 U
5688 0 0
2
44287.7 2
0
5 4071~
219 584 809 0 3 22
0 45 50 17
0
0 0 624 270
4 4071
-7 -24 21 -16
3 U3C
-6 -6 15 2
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 8 9 10 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 3 3 0
1 U
7351 0 0
2
44287.7 1
0
5 4071~
219 550 809 0 3 22
0 44 51 22
0
0 0 624 270
4 4071
-7 -24 21 -16
3 U3B
-6 -6 15 2
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 5 6 4 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 2 3 0
1 U
392 0 0
2
44287.7 0
0
4 4008
219 868 710 0 14 29
0 101 102 103 52 54 55 56 57 104
40 41 42 43 105
0
0 0 4848 782
4 4008
-14 -60 14 -52
3 U17
50 -7 71 1
0
15 DVDD=16;DGND=8;
126 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 1 3 5 7 15 2 4 6 9
10 11 12 13 14 1 3 5 7 15
2 4 6 9 10 11 12 13 14 0
65 0 0 512 0 0 0 0
1 U
5788 0 0
2
44287.7 0
0
9 Inverter~
13 901 523 0 2 22
0 64 67
0
0 0 624 782
6 74LS04
-21 -19 21 -11
4 U15E
-9 -8 19 0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 11 10 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 5 6 0
1 U
4290 0 0
2
44287.7 3
0
9 Inverter~
13 926 523 0 2 22
0 65 66
0
0 0 624 782
6 74LS04
-21 -19 21 -11
4 U15D
-9 -8 19 0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 9 8 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 4 6 0
1 U
3479 0 0
2
44287.7 2
0
9 Inverter~
13 877 523 0 2 22
0 63 68
0
0 0 624 782
6 74LS04
-21 -19 21 -11
4 U15C
-9 -8 19 0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 5 6 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 3 6 0
1 U
886 0 0
2
44287.7 1
0
9 Inverter~
13 852 523 0 2 22
0 62 69
0
0 0 624 782
6 74LS04
-21 -19 21 -11
4 U15B
-9 -8 19 0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 3 4 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 2 6 0
1 U
8133 0 0
2
44287.7 0
0
13 Quad 3-State~
48 512 588 0 9 19
0 74 75 76 77 61 60 59 58 79
0
0 0 4720 270
8 QUAD3STA
-28 -44 28 -36
3 U11
42 -1 63 7
0
15 DVCC=16;DGND=8;
85 %D [%16bi %8bi %1i %2i %3i %4i %9i]
+ [%16bo %1o %2o %3o %4o %9o %5o %6o %7o %8o] %M
0
12 type:digital
5 DIP16
19

0 1 2 3 4 5 6 7 8 9
1 2 3 4 5 6 7 8 9 0
65 0 0 0 1 0 0 0
1 U
8564 0 0
2
44287.7 0
0
13 Quad 3-State~
48 877 592 0 9 19
0 66 67 68 69 57 56 55 54 78
0
0 0 4720 270
8 QUAD3STA
-28 -44 28 -36
3 U13
42 -1 63 7
0
15 DVCC=16;DGND=8;
85 %D [%16bi %8bi %1i %2i %3i %4i %9i]
+ [%16bo %1o %2o %3o %4o %9o %5o %6o %7o %8o] %M
0
12 type:digital
5 DIP16
19

0 1 2 3 4 5 6 7 8 9
1 2 3 4 5 6 7 8 9 0
65 0 0 0 1 0 0 0
1 U
5876 0 0
2
44287.7 0
0
9 Inverter~
13 831 576 0 2 22
0 52 78
0
0 0 624 782
6 74LS04
-21 -19 21 -11
4 U15A
-9 -8 19 0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 1 6 0
1 U
6693 0 0
2
44287.7 0
0
9 Inverter~
13 459 572 0 2 22
0 53 79
0
0 0 624 782
6 74LS04
-21 -19 21 -11
3 U8F
-6 -8 15 0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 13 12 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 6 4 0
1 U
4551 0 0
2
44287.7 0
0
9 Inverter~
13 482 523 0 2 22
0 70 77
0
0 0 624 782
6 74LS04
-21 -19 21 -11
3 U8B
-6 -8 15 0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 3 4 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 2 4 0
1 U
5790 0 0
2
44287.7 3
0
9 Inverter~
13 507 523 0 2 22
0 71 76
0
0 0 624 782
6 74LS04
-21 -19 21 -11
3 U8C
-6 -8 15 0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 5 6 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 3 4 0
1 U
3845 0 0
2
44287.7 2
0
9 Inverter~
13 556 523 0 2 22
0 73 74
0
0 0 624 782
6 74LS04
-21 -19 21 -11
3 U8D
-6 -8 15 0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 9 8 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 4 4 0
1 U
8294 0 0
2
44287.7 1
0
9 Inverter~
13 531 523 0 2 22
0 72 75
0
0 0 624 782
6 74LS04
-21 -19 21 -11
3 U8E
-6 -8 15 0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 11 10 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 5 4 0
1 U
7344 0 0
2
44287.7 0
0
4 4008
219 501 705 0 14 29
0 106 107 108 53 58 59 60 61 109
48 49 50 51 110
0
0 0 4848 782
4 4008
-14 -60 14 -52
3 U10
50 -7 71 1
0
15 DVDD=16;DGND=8;
126 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 1 3 5 7 15 2 4 6 9
10 11 12 13 14 1 3 5 7 15
2 4 6 9 10 11 12 13 14 0
65 0 0 512 0 0 0 0
1 U
3552 0 0
2
44287.7 0
0
10 Buffer 3S~
219 806 255 0 3 22
0 83 80 52
0
0 0 624 270
8 BUFFER3S
-27 -51 29 -43
3 U9B
13 -5 34 3
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
0
22

0 5 4 6 2 1 3 5 4 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 5 0
1 U
5966 0 0
2
44287.7 2
0
14 Logic Display~
6 788 212 0 1 2
10 83
0
0 0 53856 0
6 100MEG
3 -16 45 -8
3 L11
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
3284 0 0
2
44287.7 0
0
14 Logic Display~
6 324 273 0 1 2
10 80
0
0 0 53856 0
6 100MEG
3 -16 45 -8
3 L10
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
570 0 0
2
44287.7 0
0
14 Logic Display~
6 513 215 0 1 2
10 84
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L9
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
3987 0 0
2
44287.7 0
0
10 Buffer 3S~
219 531 258 0 3 22
0 84 80 53
0
0 0 624 270
8 BUFFER3S
-27 -51 29 -43
3 U9A
13 -5 34 3
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
0
22

0 2 1 3 2 1 3 5 4 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 5 0
1 U
7285 0 0
2
44287.7 0
0
14 Logic Display~
6 933 219 0 1 2
10 85
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L5
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
3584 0 0
2
44287.7 7
0
14 Logic Display~
6 900 219 0 1 2
10 86
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L6
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
3181 0 0
2
44287.7 5
0
14 Logic Display~
6 866 217 0 1 2
10 87
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L7
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
3154 0 0
2
44287.7 3
0
14 Logic Display~
6 831 216 0 1 2
10 88
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L8
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
3397 0 0
2
44287.7 1
0
9 Inverter~
13 380 293 0 2 22
0 80 81
0
0 0 624 692
6 74LS04
-21 -19 21 -11
3 U8A
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 1 4 0
1 U
3654 0 0
2
44287.7 1
0
14 Logic Display~
6 663 218 0 1 2
10 97
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L4
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
6959 0 0
2
44287.7 1
0
14 Logic Display~
6 630 218 0 1 2
10 98
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L3
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
3688 0 0
2
44287.7 1
0
14 Logic Display~
6 596 216 0 1 2
10 99
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L2
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
7228 0 0
2
44287.7 1
0
14 Logic Display~
6 561 215 0 1 2
10 100
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
6996 0 0
2
44287.7 1
0
7 Pulser~
4 247 360 0 10 12
0 111 112 82 113 0 0 5 5 3
8
0
0 0 4656 0
0
2 V2
-7 -28 7 -20
0
0
0
0
0
4 SIP2
9

0 1 2 3 4 1 2 3 4 0
0 0 0 512 0 0 0 0
1 V
3550 0 0
2
44287.7 0
0
159
1 3 2 0 0 4224 0 19 20 0 0 2
363 1416
363 1417
0 2 3 0 0 4224 0 0 20 57 0 4
376 1190
376 1281
354 1281
354 1368
0 1 4 0 0 4224 0 0 20 44 0 3
610 1325
372 1325
372 1368
1 0 5 0 0 0 0 21 0 0 13 2
1216 1106
1216 1106
1 0 6 0 0 0 0 22 0 0 12 2
1176 1103
1176 1103
1 0 7 0 0 4096 0 40 0 0 9 2
1155 1217
1279 1217
3 0 8 0 0 4096 0 37 0 0 8 2
1185 1311
1185 1354
2 2 8 0 0 4224 0 40 36 0 0 3
1155 1235
1155 1354
1228 1354
0 1 7 0 0 8192 0 0 36 67 0 5
1225 980
1279 980
1279 1345
1246 1345
1246 1354
2 0 5 0 0 4096 0 39 0 0 13 2
1154 1191
1194 1191
1 0 6 0 0 4096 0 39 0 0 12 2
1154 1173
1176 1173
3 2 6 0 0 8320 0 65 37 0 0 4
654 839
654 919
1176 919
1176 1262
1 3 5 0 0 4224 0 37 57 0 0 4
1194 1262
1194 1117
1216 1117
1216 1059
1 3 9 0 0 4224 0 23 36 0 0 2
1237 1402
1237 1403
1 0 10 0 0 4096 0 24 0 0 26 2
1005 1104
1004 1104
1 0 11 0 0 0 0 25 0 0 25 2
986 1105
986 1105
1 0 12 0 0 12416 0 41 0 0 20 4
1056 1349
1056 1319
1023 1319
1023 1209
1 0 12 0 0 0 0 26 0 0 20 2
1036 1202
1036 1201
1 3 13 0 0 4224 0 27 41 0 0 2
1047 1397
1047 1398
3 1 12 0 0 0 0 38 45 0 0 4
1040 1201
1023 1201
1023 1212
953 1212
2 0 14 0 0 4224 0 45 0 0 22 3
953 1230
953 1348
995 1348
3 2 14 0 0 0 0 42 41 0 0 3
995 1306
995 1349
1038 1349
2 0 10 0 0 4096 0 44 0 0 26 2
951 1186
1004 1186
1 0 11 0 0 4096 0 44 0 0 25 2
951 1168
986 1168
3 2 11 0 0 8320 0 66 42 0 0 6
620 839
620 931
914 931
914 1076
986 1076
986 1257
3 1 10 0 0 8320 0 58 42 0 0 3
991 1059
1004 1059
1004 1257
1 0 15 0 0 0 0 28 0 0 32 2
841 1196
841 1196
1 0 16 0 0 4096 0 30 0 0 38 2
791 1106
789 1106
1 0 17 0 0 4096 0 31 0 0 37 2
768 1106
771 1106
1 3 18 0 0 4224 0 29 50 0 0 2
832 1400
832 1396
1 0 15 0 0 4096 0 46 0 0 32 2
734 1211
841 1211
1 3 15 0 0 4224 0 50 43 0 0 3
841 1347
841 1196
850 1196
0 2 19 0 0 8320 0 0 46 34 0 3
780 1347
734 1347
734 1229
2 3 19 0 0 0 0 50 49 0 0 3
823 1347
780 1347
780 1304
2 0 16 0 0 4096 0 47 0 0 38 2
736 1184
789 1184
1 0 17 0 0 4096 0 47 0 0 37 2
736 1166
771 1166
3 2 17 0 0 12416 0 67 49 0 0 4
587 839
587 939
771 939
771 1255
1 3 16 0 0 4224 0 49 59 0 0 4
789 1255
789 1073
799 1073
799 1060
1 3 20 0 0 4224 0 34 56 0 0 2
601 1400
601 1396
1 0 21 0 0 0 0 32 0 0 50 2
594 1104
594 1104
1 0 22 0 0 4096 0 33 0 0 49 2
537 1106
538 1106
1 0 4 0 0 0 0 35 0 0 43 2
621 1194
621 1194
3 0 4 0 0 0 0 48 0 0 44 3
632 1194
609 1194
609 1206
1 1 4 0 0 0 0 53 56 0 0 3
516 1206
610 1206
610 1347
3 0 23 0 0 4096 0 55 0 0 46 2
547 1308
547 1347
2 2 23 0 0 8320 0 53 56 0 0 4
516 1224
524 1224
524 1347
592 1347
2 0 21 0 0 4096 0 52 0 0 50 2
515 1180
556 1180
1 0 22 0 0 4096 0 52 0 0 49 2
515 1162
538 1162
3 2 22 0 0 4224 0 68 55 0 0 4
553 839
553 1098
538 1098
538 1259
1 3 21 0 0 4224 0 55 60 0 0 4
556 1259
556 1121
594 1121
594 1058
2 3 24 0 0 8320 0 38 40 0 0 4
1086 1210
1101 1210
1101 1226
1110 1226
3 1 25 0 0 12416 0 39 38 0 0 4
1109 1182
1101 1182
1101 1192
1086 1192
2 3 26 0 0 8320 0 43 45 0 0 3
896 1205
908 1205
908 1221
3 1 27 0 0 4224 0 44 43 0 0 3
906 1177
906 1187
896 1187
2 3 28 0 0 8320 0 48 46 0 0 3
678 1203
689 1203
689 1220
3 1 29 0 0 8320 0 47 48 0 0 3
691 1175
691 1185
678 1185
1 3 3 0 0 0 0 54 51 0 0 3
376 1181
376 1190
401 1190
2 3 30 0 0 8320 0 51 53 0 0 4
447 1199
462 1199
462 1215
471 1215
3 1 31 0 0 12416 0 52 51 0 0 4
470 1171
462 1171
462 1181
447 1181
3 2 32 0 0 8320 0 64 60 0 0 4
934 859
934 954
585 954
585 1009
2 3 33 0 0 8320 0 59 63 0 0 4
790 1011
790 967
968 967
968 859
2 3 34 0 0 12416 0 58 62 0 0 4
982 1010
982 968
1001 968
1001 859
2 3 35 0 0 8320 0 57 61 0 0 4
1207 1010
1207 968
1035 968
1035 859
1 0 7 0 0 0 0 1 0 0 67 4
334 921
378 921
378 980
604 980
1 0 7 0 0 0 0 58 0 0 67 2
1000 1010
1000 980
1 0 7 0 0 0 0 59 0 0 67 2
808 1011
808 980
1 1 7 0 0 8320 0 57 60 0 0 4
1225 1010
1225 980
603 980
603 1009
1 8 36 0 0 12416 0 64 13 0 0 4
943 813
943 729
1028 729
1028 617
1 7 37 0 0 12416 0 63 13 0 0 4
977 813
977 739
1040 739
1040 617
1 6 38 0 0 12416 0 62 13 0 0 4
1010 813
1010 747
1052 747
1052 617
1 5 39 0 0 12416 0 61 13 0 0 4
1044 813
1044 756
1064 756
1064 617
10 2 40 0 0 8320 0 69 61 0 0 4
879 740
879 764
1026 764
1026 813
2 11 41 0 0 8320 0 62 69 0 0 4
992 813
992 771
870 771
870 740
12 2 42 0 0 8320 0 69 63 0 0 4
861 740
861 784
959 784
959 813
13 2 43 0 0 8320 0 69 64 0 0 4
852 740
852 798
925 798
925 813
8 1 44 0 0 12416 0 14 68 0 0 6
646 614
646 666
584 666
584 741
562 741
562 793
1 7 45 0 0 4224 0 67 14 0 0 4
596 793
596 683
658 683
658 614
1 6 46 0 0 4224 0 66 14 0 0 4
629 793
629 693
670 693
670 614
1 5 47 0 0 12416 0 65 14 0 0 4
663 793
663 709
682 709
682 614
10 2 48 0 0 8320 0 82 65 0 0 4
512 735
512 751
645 751
645 793
2 11 49 0 0 8320 0 66 82 0 0 4
611 793
611 760
503 760
503 735
12 2 50 0 0 8320 0 82 67 0 0 4
494 735
494 770
578 770
578 793
2 13 51 0 0 8320 0 68 82 0 0 4
544 793
544 782
485 782
485 735
4 0 52 0 0 12288 0 69 0 0 107 4
861 676
861 642
805 642
805 543
0 4 53 0 0 8192 0 0 82 117 0 5
462 540
426 540
426 659
494 659
494 671
5 8 54 0 0 4224 0 69 75 0 0 4
870 676
870 641
874 641
874 619
6 7 55 0 0 4224 0 69 75 0 0 4
879 676
879 646
886 646
886 619
7 6 56 0 0 12416 0 69 75 0 0 4
888 676
888 654
898 654
898 619
8 5 57 0 0 12416 0 69 75 0 0 4
897 676
897 665
910 665
910 619
5 8 58 0 0 4224 0 82 74 0 0 4
503 671
503 629
509 629
509 615
6 7 59 0 0 4224 0 82 74 0 0 4
512 671
512 637
521 637
521 615
7 6 60 0 0 12416 0 82 74 0 0 4
521 671
521 644
533 644
533 615
8 5 61 0 0 12416 0 82 74 0 0 4
530 671
530 649
545 649
545 615
0 4 62 0 0 4224 0 0 13 101 0 3
855 484
1028 484
1028 569
0 3 63 0 0 4224 0 0 13 100 0 3
880 478
1040 478
1040 569
0 2 64 0 0 4224 0 0 13 99 0 3
904 472
1052 472
1052 569
0 1 65 0 0 4224 0 0 13 98 0 3
929 465
1064 465
1064 569
1 5 65 0 0 0 0 71 15 0 0 3
929 505
929 428
916 428
1 6 64 0 0 0 0 70 15 0 0 2
904 505
904 428
1 7 63 0 0 0 0 72 15 0 0 4
880 505
880 466
892 466
892 428
1 8 62 0 0 0 0 73 15 0 0 4
855 505
855 458
880 458
880 428
0 9 52 0 0 4096 0 0 13 107 0 3
805 494
992 494
992 593
1 2 66 0 0 8320 0 75 71 0 0 3
910 571
929 571
929 541
2 2 67 0 0 12416 0 75 70 0 0 4
898 571
898 558
904 558
904 541
3 2 68 0 0 4224 0 75 72 0 0 4
886 571
886 554
880 554
880 541
2 4 69 0 0 4224 0 73 75 0 0 4
855 541
855 560
874 560
874 571
3 1 52 0 0 4224 0 83 76 0 0 4
805 271
805 545
834 545
834 558
0 9 53 0 0 8320 0 0 14 117 0 4
530 427
588 427
588 590
610 590
4 0 70 0 0 12288 0 14 0 0 116 4
646 566
646 552
621 552
621 456
3 0 71 0 0 12288 0 14 0 0 115 4
658 566
658 537
633 537
633 464
2 0 72 0 0 12288 0 14 0 0 114 4
670 566
670 524
643 524
643 471
1 0 73 0 0 4096 0 14 0 0 113 4
682 566
682 511
656 511
656 483
1 5 73 0 0 8320 0 80 16 0 0 4
559 505
559 483
657 483
657 433
1 6 72 0 0 8320 0 81 16 0 0 4
534 505
534 471
645 471
645 433
1 7 71 0 0 8320 0 79 16 0 0 4
510 505
510 464
633 464
633 433
1 8 70 0 0 8320 0 78 16 0 0 4
485 505
485 456
621 456
621 433
3 1 53 0 0 0 0 87 77 0 0 4
530 274
530 427
462 427
462 554
1 2 74 0 0 8320 0 74 80 0 0 3
545 567
559 567
559 541
2 2 75 0 0 8320 0 74 81 0 0 3
533 567
534 567
534 541
2 3 76 0 0 8320 0 79 74 0 0 3
510 541
521 541
521 567
2 4 77 0 0 8320 0 78 74 0 0 4
485 541
485 559
509 559
509 567
2 9 78 0 0 8320 0 76 75 0 0 3
834 594
834 595
838 595
2 9 79 0 0 8320 0 77 74 0 0 3
462 590
462 591
473 591
0 2 80 0 0 8192 0 0 87 146 0 3
348 293
348 259
519 259
0 2 80 0 0 8320 0 0 83 146 0 5
335 293
335 347
777 347
777 256
794 256
0 9 81 0 0 8320 0 0 17 127 0 5
563 308
563 340
832 340
832 304
844 304
2 9 81 0 0 0 0 92 18 0 0 4
401 293
488 293
488 308
585 308
0 9 82 0 0 8320 0 0 15 147 0 5
571 409
571 372
832 372
832 404
850 404
0 1 83 0 0 4224 0 0 84 130 0 3
805 234
788 234
788 230
1 1 83 0 0 0 0 83 2 0 0 2
805 241
805 226
1 0 80 0 0 0 0 85 0 0 146 2
324 291
324 293
0 1 84 0 0 4224 0 0 86 133 0 3
530 237
513 237
513 233
1 1 84 0 0 0 0 87 3 0 0 2
530 244
530 229
1 0 85 0 0 8320 0 17 0 0 142 3
916 280
939 280
939 246
2 0 86 0 0 12416 0 17 0 0 143 4
904 280
904 273
907 273
907 246
3 0 87 0 0 12416 0 17 0 0 144 4
892 280
892 274
875 274
875 244
4 0 88 0 0 4224 0 17 0 0 145 3
880 280
840 280
840 243
4 8 89 0 0 4224 0 15 17 0 0 2
880 380
880 328
3 7 90 0 0 4224 0 15 17 0 0 2
892 380
892 328
2 6 91 0 0 4224 0 15 17 0 0 2
904 380
904 328
1 5 92 0 0 4224 0 15 17 0 0 2
916 380
916 328
1 1 85 0 0 0 0 4 88 0 0 4
950 233
950 246
933 246
933 237
1 1 86 0 0 0 0 5 89 0 0 4
917 233
917 246
900 246
900 237
1 1 87 0 0 0 0 6 90 0 0 4
883 231
883 244
866 244
866 235
1 1 88 0 0 0 0 7 91 0 0 4
848 230
848 243
831 243
831 234
1 1 80 0 0 0 0 92 8 0 0 2
365 293
314 293
3 9 82 0 0 0 0 97 16 0 0 4
271 351
413 351
413 409
591 409
4 8 93 0 0 4224 0 16 18 0 0 2
621 385
621 332
3 7 94 0 0 4224 0 16 18 0 0 2
633 385
633 332
2 6 95 0 0 4224 0 16 18 0 0 2
645 385
645 332
1 5 96 0 0 4224 0 16 18 0 0 2
657 385
657 332
1 0 97 0 0 12416 0 18 0 0 156 4
657 284
657 265
671 265
671 245
2 0 98 0 0 12416 0 18 0 0 157 4
645 284
645 269
640 269
640 245
3 0 99 0 0 12416 0 18 0 0 158 4
633 284
633 273
605 273
605 243
4 0 100 0 0 4224 0 18 0 0 159 3
621 284
569 284
569 242
1 1 97 0 0 0 0 9 93 0 0 4
680 232
680 245
663 245
663 236
1 1 98 0 0 0 0 10 94 0 0 4
647 232
647 245
630 245
630 236
1 1 99 0 0 0 0 11 95 0 0 4
613 230
613 243
596 243
596 234
1 1 100 0 0 0 0 12 96 0 0 4
578 229
578 242
561 242
561 233
4
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 31
201 1406 350 1450
211 1414 339 1446
31 Vai ser Overflow 
se der 1 =>
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 21
250 1108 439 1132
260 1116 428 1132
21 Vai 1(Fora do numero)
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 12
465 1399 582 1423
475 1407 571 1423
12 Resultado =>
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 31
244 831 353 895
254 839 342 887
31 Controle
0 - Soma
1 - Subtrai
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0

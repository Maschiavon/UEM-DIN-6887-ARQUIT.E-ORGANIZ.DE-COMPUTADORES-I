CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 1 100 10
176 80 1918 1019
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
0 4 0.500000 0.500000
344 176 457 273
42991634 0
0
6 Title:
5 Name:
0
0
0
44
13 Logic Switch~
5 267 282 0 10 11
0 30 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V5
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
634 0 0
2
44287.8 0
0
13 Logic Switch~
5 250 239 0 10 11
0 32 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V3
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
8956 0 0
2
44287.8 0
0
13 Logic Switch~
5 121 283 0 10 11
0 33 0 0 0 0 0 0 0 0
1
0
0 0 21360 270
2 5V
-6 -21 8 -13
2 V1
-6 -31 8 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
3342 0 0
2
44287.8 0
0
13 Logic Switch~
5 75 284 0 10 11
0 34 0 0 0 0 0 0 0 0
1
0
0 0 21360 270
2 5V
-6 -21 8 -13
2 V4
-6 -31 8 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
3549 0 0
2
44287.8 0
0
14 Logic Display~
6 926 213 0 1 2
10 13
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 F4
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
9177 0 0
2
44287.8 2
0
14 Logic Display~
6 1014 207 0 1 2
10 12
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 F5
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
3387 0 0
2
44287.8 1
0
14 Logic Display~
6 1107 210 0 1 2
10 11
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 F6
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
351 0 0
2
44287.8 0
0
14 Logic Display~
6 760 220 0 1 2
10 15
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 F2
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
3127 0 0
2
44287.8 2
0
9 8-In NOR~
219 755 315 0 9 19
0 8 5 4 37 38 39 40 41 16
0
0 0 624 90
4 4078
-7 -24 21 -16
2 U9
9 -8 23 0
0
15 DVDD=14;DGND=7;
97 %D [%14bi %7bi %1i %2i %3i %4i %5i %6i %7i %8i]
+ [%14bo %1o %2o %3o %4o %5o %6o %7o %8o %9o] %M
0
12 type:digital
5 DIP14
19

0 2 3 4 5 9 10 11 12 13
2 3 4 5 9 10 11 12 13 0
65 0 0 512 0 0 0 0
1 U
559 0 0
2
44287.8 1
0
9 Inverter~
13 757 255 0 2 22
0 16 15
0
0 0 624 90
6 74LS04
-21 -19 21 -11
3 U6F
16 -2 37 6
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 13 12 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 6 3 0
1 U
8488 0 0
2
44287.8 0
0
9 Inverter~
13 1106 253 0 2 22
0 17 11
0
0 0 624 90
6 74LS04
-21 -19 21 -11
4 U11D
13 -2 41 6
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 9 8 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 4 6 0
1 U
3392 0 0
2
44287.8 1
0
9 8-In NOR~
219 1104 313 0 9 19
0 9 7 5 3 42 43 44 45 17
0
0 0 624 90
4 4078
-7 -24 21 -16
3 U14
6 -8 27 0
0
15 DVDD=14;DGND=7;
97 %D [%14bi %7bi %1i %2i %3i %4i %5i %6i %7i %8i]
+ [%14bo %1o %2o %3o %4o %5o %6o %7o %8o %9o] %M
0
12 type:digital
5 DIP14
19

0 2 3 4 5 9 10 11 12 13
2 3 4 5 9 10 11 12 13 0
65 0 0 512 0 0 0 0
1 U
3952 0 0
2
44287.8 0
0
9 Inverter~
13 1011 254 0 2 22
0 18 12
0
0 0 624 90
6 74LS04
-21 -19 21 -11
4 U11C
13 -2 41 6
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 5 6 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 3 6 0
1 U
8186 0 0
2
44287.8 1
0
9 8-In NOR~
219 1009 314 0 9 19
0 9 6 3 46 47 48 49 50 18
0
0 0 624 90
4 4078
-7 -24 21 -16
3 U13
6 -8 27 0
0
15 DVDD=14;DGND=7;
97 %D [%14bi %7bi %1i %2i %3i %4i %5i %6i %7i %8i]
+ [%14bo %1o %2o %3o %4o %5o %6o %7o %8o %9o] %M
0
12 type:digital
5 DIP14
19

0 2 3 4 5 9 10 11 12 13
2 3 4 5 9 10 11 12 13 0
65 0 0 512 0 0 0 0
1 U
6571 0 0
2
44287.8 0
0
9 Inverter~
13 926 255 0 2 22
0 19 13
0
0 0 624 90
6 74LS04
-21 -19 21 -11
4 U11B
13 -2 41 6
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 3 4 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 2 6 0
1 U
6167 0 0
2
44287.8 1
0
9 8-In NOR~
219 924 315 0 9 19
0 8 3 51 52 53 54 55 56 19
0
0 0 624 90
4 4078
-7 -24 21 -16
3 U12
6 -8 27 0
0
15 DVDD=14;DGND=7;
97 %D [%14bi %7bi %1i %2i %3i %4i %5i %6i %7i %8i]
+ [%14bo %1o %2o %3o %4o %5o %6o %7o %8o %9o] %M
0
12 type:digital
5 DIP14
19

0 2 3 4 5 9 10 11 12 13
2 3 4 5 9 10 11 12 13 0
65 0 0 512 0 0 0 0
1 U
3566 0 0
2
44287.8 0
0
9 Inverter~
13 840 250 0 2 22
0 20 14
0
0 0 624 90
6 74LS04
-21 -19 21 -11
4 U11A
13 -2 41 6
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 1 6 0
1 U
3371 0 0
2
44287.8 1
0
9 8-In NOR~
219 838 310 0 9 19
0 10 7 5 4 57 58 59 60 20
0
0 0 624 90
4 4078
-7 -24 21 -16
3 U10
6 -8 27 0
0
15 DVDD=14;DGND=7;
97 %D [%14bi %7bi %1i %2i %3i %4i %5i %6i %7i %8i]
+ [%14bo %1o %2o %3o %4o %5o %6o %7o %8o %9o] %M
0
12 type:digital
5 DIP14
19

0 2 3 4 5 9 10 11 12 13
2 3 4 5 9 10 11 12 13 0
65 0 0 512 0 0 0 0
1 U
4395 0 0
2
44287.8 0
0
14 Logic Display~
6 843 215 0 1 2
10 14
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 F3
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
6822 0 0
2
44287.8 0
0
14 Logic Display~
6 678 216 0 1 2
10 21
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 F1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
8953 0 0
2
44287.8 2
0
9 8-In NOR~
219 671 314 0 9 19
0 10 6 4 61 62 63 64 65 22
0
0 0 624 90
4 4078
-7 -24 21 -16
2 U8
9 -8 23 0
0
15 DVDD=14;DGND=7;
97 %D [%14bi %7bi %1i %2i %3i %4i %5i %6i %7i %8i]
+ [%14bo %1o %2o %3o %4o %5o %6o %7o %8o %9o] %M
0
12 type:digital
5 DIP14
19

0 2 3 4 5 9 10 11 12 13
2 3 4 5 9 10 11 12 13 0
65 0 0 512 0 0 0 0
1 U
4635 0 0
2
44287.8 1
0
9 Inverter~
13 673 254 0 2 22
0 22 21
0
0 0 624 90
6 74LS04
-21 -19 21 -11
3 U6E
16 -2 37 6
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 11 10 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 5 3 0
1 U
6596 0 0
2
44287.8 0
0
9 2-In AND~
219 466 543 0 3 22
0 25 2 6
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U7D
-13 -11 8 -3
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 5 0
1 U
3813 0 0
2
44287.8 3
0
9 2-In AND~
219 467 580 0 3 22
0 25 23 5
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U7C
-13 -14 8 -6
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 5 0
1 U
5639 0 0
2
44287.8 2
0
9 2-In AND~
219 468 619 0 3 22
0 24 2 4
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U7B
-13 -14 8 -6
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 5 0
1 U
429 0 0
2
44287.8 1
0
9 2-In AND~
219 466 657 0 3 22
0 24 23 3
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U7A
-13 -14 8 -6
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 5 0
1 U
5832 0 0
2
44287.8 0
0
9 2-In AND~
219 467 501 0 3 22
0 26 23 7
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U4D
-13 -14 8 -6
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 4 0
1 U
8856 0 0
2
44287.8 0
0
9 2-In AND~
219 469 463 0 3 22
0 26 2 8
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U4C
-13 -14 8 -6
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 4 0
1 U
469 0 0
2
44287.8 0
0
9 2-In AND~
219 468 424 0 3 22
0 27 23 9
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U4B
-13 -14 8 -6
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 4 0
1 U
4529 0 0
2
44287.8 0
0
9 2-In AND~
219 467 387 0 3 22
0 27 2 10
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U4A
-13 -11 8 -3
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 4 0
1 U
88 0 0
2
44287.8 0
0
9 Inverter~
13 389 337 0 2 22
0 23 2
0
0 0 624 270
6 74LS04
-21 -19 21 -11
3 U6D
16 -8 37 0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 9 8 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 4 3 0
1 U
3894 0 0
2
44287.8 0
0
14 Logic Display~
6 332 170 0 1 2
10 29
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L5
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
6890 0 0
2
44287.8 0
0
9 2-In AND~
219 201 395 0 3 22
0 36 35 27
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U5A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 2 0
1 U
3257 0 0
2
44287.8 3
0
9 2-In AND~
219 203 444 0 3 22
0 36 33 26
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U5B
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 2 0
1 U
6612 0 0
2
44287.8 2
0
9 2-In AND~
219 204 492 0 3 22
0 34 35 25
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U5C
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 2 0
1 U
3556 0 0
2
44287.8 1
0
9 2-In AND~
219 206 542 0 3 22
0 34 33 24
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U5D
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 2 0
1 U
9143 0 0
2
44287.8 0
0
9 Inverter~
13 125 341 0 2 22
0 33 35
0
0 0 624 270
6 74LS04
-21 -19 21 -11
3 U6B
-7 -9 14 -1
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 3 4 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 2 3 0
1 U
8186 0 0
2
44287.8 0
0
9 Inverter~
13 56 342 0 2 22
0 34 36
0
0 0 624 270
6 74LS04
-21 -19 21 -11
3 U6A
-6 -14 15 -6
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 1 3 0
1 U
3754 0 0
2
44287.8 0
0
14 Logic Display~
6 142 278 0 1 2
10 33
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L3
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
8708 0 0
2
44287.8 0
0
14 Logic Display~
6 55 278 0 1 2
10 34
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L2
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
3338 0 0
2
44287.8 0
0
10 Buffer 3S~
219 370 191 0 3 22
0 29 32 23
0
0 0 624 0
8 BUFFER3S
-27 -51 29 -43
3 U1B
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
0
22

0 5 4 6 2 1 3 5 4 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 1 0
1 U
5546 0 0
2
44287.8 0
0
12 D Flip-Flop~
219 291 227 0 4 9
0 31 28 66 29
0
0 0 4720 0
3 DFF
-10 -53 11 -45
2 U3
-7 -55 7 -47
0
14 DVCC=6;DGND=5;
47 %D [%6bi %5bi %1i %2i][%6bo %1o %2o %3o %4o] %M
0
11 typeDigital
4 DIP6
9

0 1 2 3 4 1 2 3 4 0
65 0 0 512 1 0 0 0
1 U
3295 0 0
2
44287.8 0
0
4 4008
219 496 259 0 14 29
0 67 68 69 29 70 71 72 30 73
31 74 75 76 77
0
0 0 4848 0
4 4008
-14 -60 14 -52
2 U2
-7 -61 7 -53
0
15 DVDD=16;DGND=8;
126 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 1 3 5 7 15 2 4 6 9
10 11 12 13 14 1 3 5 7 15
2 4 6 9 10 11 12 13 14 0
65 0 0 512 0 0 0 0
1 U
4923 0 0
2
44287.8 0
0
7 Pulser~
4 63 171 0 10 12
0 78 79 28 80 0 0 5 5 3
7
0
0 0 4656 0
0
2 V2
-7 -28 7 -20
0
0
0
0
0
4 SIP2
9

0 1 2 3 4 1 2 3 4 0
0 0 0 512 0 0 0 0
1 V
3248 0 0
2
44287.8 0
0
68
0 2 2 0 0 4096 0 0 25 37 0 3
396 552
396 628
444 628
0 4 3 0 0 8192 0 0 12 3 0 3
1002 657
1106 657
1106 336
0 3 3 0 0 0 0 0 14 4 0 3
907 657
1002 657
1002 337
3 2 3 0 0 4224 0 26 16 0 0 3
487 657
908 657
908 338
0 4 4 0 0 8336 0 0 18 6 0 3
748 619
840 619
840 333
0 3 4 0 0 0 0 0 9 7 0 3
662 619
748 619
748 338
3 3 4 0 0 0 0 25 21 0 0 3
489 619
664 619
664 337
0 3 5 0 0 4224 0 0 12 9 0 3
830 580
1097 580
1097 336
0 3 5 0 0 0 0 0 18 10 0 3
738 580
831 580
831 333
3 2 5 0 0 0 0 24 9 0 0 3
488 580
739 580
739 338
0 2 6 0 0 4224 0 0 14 12 0 3
655 543
993 543
993 337
3 2 6 0 0 0 0 23 21 0 0 3
487 543
655 543
655 337
2 0 7 0 0 8192 0 12 0 0 14 3
1088 336
1088 501
822 501
3 2 7 0 0 4224 0 27 18 0 0 3
488 501
822 501
822 333
1 0 8 0 0 8192 0 16 0 0 16 3
899 338
899 463
730 463
3 1 8 0 0 4224 0 28 9 0 0 3
490 463
730 463
730 338
0 1 9 0 0 4096 0 0 12 18 0 3
984 424
1079 424
1079 336
3 1 9 0 0 4224 0 29 14 0 0 3
489 424
984 424
984 337
0 1 10 0 0 4224 0 0 18 20 0 3
646 387
813 387
813 333
3 1 10 0 0 0 0 30 21 0 0 3
488 387
646 387
646 337
1 2 11 0 0 4224 0 7 11 0 0 4
1107 228
1107 236
1109 236
1109 235
1 2 12 0 0 4224 0 6 13 0 0 4
1014 225
1014 237
1014 237
1014 236
1 2 13 0 0 4224 0 5 15 0 0 3
926 231
926 237
929 237
1 2 14 0 0 4224 0 19 17 0 0 2
843 233
843 232
2 1 15 0 0 4224 0 10 8 0 0 2
760 237
760 238
1 9 16 0 0 4224 0 10 9 0 0 4
760 273
760 283
761 283
761 282
1 9 17 0 0 4224 0 11 12 0 0 4
1109 271
1109 281
1110 281
1110 280
1 9 18 0 0 4224 0 13 14 0 0 4
1014 272
1014 282
1015 282
1015 281
1 9 19 0 0 4224 0 15 16 0 0 4
929 273
929 283
930 283
930 282
1 9 20 0 0 4224 0 17 18 0 0 4
843 268
843 278
844 278
844 277
1 2 21 0 0 4224 0 20 22 0 0 3
678 234
678 236
676 236
1 9 22 0 0 4224 0 22 21 0 0 4
676 272
676 282
677 282
677 281
0 2 23 0 0 4096 0 0 26 34 0 3
380 589
380 666
442 666
0 2 23 0 0 4096 0 0 24 35 0 3
380 508
380 589
443 589
0 2 23 0 0 0 0 0 27 36 0 3
380 433
380 510
443 510
0 2 23 0 0 8320 0 0 29 48 0 4
392 305
368 305
368 433
444 433
2 0 2 0 0 8320 0 23 0 0 38 3
442 552
395 552
395 472
2 0 2 0 0 0 0 28 0 0 39 3
445 472
393 472
393 396
2 2 2 0 0 0 0 30 31 0 0 3
443 396
392 396
392 355
1 0 24 0 0 4096 0 26 0 0 41 3
442 648
278 648
278 610
3 1 24 0 0 12416 0 36 25 0 0 4
227 542
278 542
278 610
444 610
1 0 25 0 0 4096 0 24 0 0 43 3
443 571
337 571
337 529
1 3 25 0 0 12416 0 23 35 0 0 4
442 534
337 534
337 492
225 492
1 0 26 0 0 4096 0 27 0 0 45 3
443 492
356 492
356 454
1 3 26 0 0 4224 0 28 34 0 0 3
445 454
224 454
224 444
1 0 27 0 0 4224 0 29 0 0 47 3
444 415
262 415
262 395
3 1 27 0 0 0 0 33 30 0 0 4
222 395
292 395
292 378
443 378
1 3 23 0 0 0 0 31 41 0 0 3
392 319
392 191
385 191
2 0 28 0 0 8192 0 42 0 0 52 3
267 209
247 209
247 162
0 4 29 0 0 8320 0 0 43 68 0 3
347 191
347 250
464 250
8 1 30 0 0 4224 0 43 1 0 0 4
464 286
284 286
284 282
279 282
3 0 28 0 0 4224 0 44 0 0 0 2
87 162
252 162
10 1 31 0 0 12416 0 43 42 0 0 8
528 268
553 268
553 129
227 129
227 194
261 194
261 191
267 191
1 0 29 0 0 0 0 32 0 0 68 2
332 188
332 191
1 2 32 0 0 8320 0 2 41 0 0 5
262 239
262 233
377 233
377 202
370 202
0 2 33 0 0 4096 0 0 36 60 0 3
147 453
147 551
182 551
0 1 34 0 0 8192 0 0 36 59 0 3
78 483
78 533
182 533
0 2 35 0 0 4224 0 0 35 62 0 3
128 404
128 501
180 501
0 1 34 0 0 8320 0 0 35 65 0 4
59 315
78 315
78 483
180 483
0 2 33 0 0 8320 0 0 34 64 0 4
128 316
147 316
147 453
179 453
1 0 36 0 0 4224 0 34 0 0 63 3
179 435
59 435
59 386
2 2 35 0 0 0 0 37 33 0 0 3
128 359
128 404
177 404
2 1 36 0 0 0 0 38 33 0 0 3
59 360
59 386
177 386
1 0 33 0 0 0 0 37 0 0 66 2
128 323
128 296
1 0 34 0 0 0 0 38 0 0 67 2
59 324
59 296
1 1 33 0 0 0 0 39 3 0 0 3
142 296
121 296
121 295
1 1 34 0 0 0 0 40 4 0 0 2
55 296
75 296
1 4 29 0 0 0 0 41 42 0 0 2
355 191
315 191
1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 18
662 136 827 160
672 144 816 160
18 F s�o as opera��es
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0

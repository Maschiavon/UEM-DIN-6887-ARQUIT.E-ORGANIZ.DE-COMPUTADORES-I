CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
1020 390 1 100 10
417 443 1183 1426
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
2 4 0.500000 0.500000
585 539 698 636
42991634 0
0
6 Title:
5 Name:
0
0
0
390
13 Logic Switch~
5 842 1587 0 10 11
0 126 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-5 -16 9 -8
3 V74
-9 -26 12 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
6230 0 0
2
5.89983e-315 0
0
13 Logic Switch~
5 830 1051 0 10 11
0 129 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-5 -16 9 -8
3 V73
-9 -26 12 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
8443 0 0
2
5.89983e-315 5.26354e-315
0
13 Logic Switch~
5 808 674 0 10 11
0 132 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-5 -16 9 -8
3 V72
-9 -26 12 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
5621 0 0
2
5.89983e-315 5.30499e-315
0
13 Logic Switch~
5 794 276 0 10 11
0 135 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-5 -16 9 -8
3 V71
-9 -26 12 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
4421 0 0
2
5.89983e-315 5.32571e-315
0
13 Logic Switch~
5 2774 1367 0 10 11
0 258 0 0 0 0 0 0 0 0
1
0
0 0 21360 270
2 5V
-6 -21 8 -13
3 V62
-9 -31 12 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
5573 0 0
2
5.89983e-315 5.34643e-315
0
13 Logic Switch~
5 2741 1367 0 10 11
0 257 0 0 0 0 0 0 0 0
1
0
0 0 21360 270
2 5V
-6 -21 8 -13
3 V63
-9 -31 12 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
8401 0 0
2
5.89983e-315 5.3568e-315
0
13 Logic Switch~
5 2710 1367 0 1 11
0 256
0
0 0 21360 270
2 0V
-6 -21 8 -13
3 V64
-9 -31 12 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
7726 0 0
2
5.89983e-315 5.36716e-315
0
13 Logic Switch~
5 2675 1367 0 10 11
0 255 0 0 0 0 0 0 0 0
1
0
0 0 21360 270
2 5V
-6 -21 8 -13
3 V65
-9 -31 12 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
9761 0 0
2
5.89983e-315 5.37752e-315
0
13 Logic Switch~
5 2388 1375 0 10 11
0 263 0 0 0 0 0 0 0 0
1
0
0 0 21360 270
2 5V
-6 -21 8 -13
3 V66
-9 -31 12 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
5847 0 0
2
5.89983e-315 5.38788e-315
0
13 Logic Switch~
5 2423 1375 0 10 11
0 264 0 0 0 0 0 0 0 0
1
0
0 0 21360 270
2 5V
-6 -21 8 -13
3 V67
-9 -31 12 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
3453 0 0
2
5.89983e-315 5.39306e-315
0
13 Logic Switch~
5 2454 1375 0 10 11
0 265 0 0 0 0 0 0 0 0
1
0
0 0 21360 270
2 5V
-6 -21 8 -13
3 V68
-9 -31 12 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
8186 0 0
2
5.89983e-315 5.39824e-315
0
13 Logic Switch~
5 2487 1375 0 10 11
0 266 0 0 0 0 0 0 0 0
1
0
0 0 21360 270
2 5V
-6 -21 8 -13
3 V69
-9 -31 12 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
4411 0 0
2
5.89983e-315 5.40342e-315
0
13 Logic Switch~
5 2763 420 0 10 11
0 274 0 0 0 0 0 0 0 0
1
0
0 0 21360 270
2 5V
-6 -21 8 -13
3 V14
-9 -31 12 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
635 0 0
2
5.89983e-315 5.4086e-315
0
13 Logic Switch~
5 2730 420 0 10 11
0 273 0 0 0 0 0 0 0 0
1
0
0 0 21360 270
2 5V
-6 -21 8 -13
3 V15
-9 -31 12 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
9584 0 0
2
5.89983e-315 5.41378e-315
0
13 Logic Switch~
5 2699 420 0 1 11
0 272
0
0 0 21360 270
2 0V
-6 -21 8 -13
3 V16
-9 -31 12 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
4959 0 0
2
5.89983e-315 5.41896e-315
0
13 Logic Switch~
5 2664 420 0 1 11
0 271
0
0 0 21360 270
2 0V
-6 -21 8 -13
3 V17
-9 -31 12 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3596 0 0
2
5.89983e-315 5.42414e-315
0
13 Logic Switch~
5 2377 428 0 1 11
0 279
0
0 0 21360 270
2 0V
-6 -21 8 -13
3 V18
-9 -31 12 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
5196 0 0
2
5.89983e-315 5.42933e-315
0
13 Logic Switch~
5 2412 428 0 10 11
0 280 0 0 0 0 0 0 0 0
1
0
0 0 21360 270
2 5V
-6 -21 8 -13
3 V19
-9 -31 12 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3372 0 0
2
5.89983e-315 5.43192e-315
0
13 Logic Switch~
5 2443 428 0 10 11
0 281 0 0 0 0 0 0 0 0
1
0
0 0 21360 270
2 5V
-6 -21 8 -13
3 V20
-9 -31 12 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
6254 0 0
2
5.89983e-315 5.43451e-315
0
13 Logic Switch~
5 2476 428 0 1 11
0 282
0
0 0 21360 270
2 0V
-6 -21 8 -13
3 V21
-9 -31 12 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
6163 0 0
2
5.89983e-315 5.4371e-315
0
13 Logic Switch~
5 2778 1680 0 10 11
0 322 0 0 0 0 0 0 0 0
1
0
0 0 21360 270
2 5V
-6 -21 8 -13
3 V61
-9 -31 12 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
4439 0 0
2
5.89983e-315 5.43969e-315
0
13 Logic Switch~
5 2745 1680 0 10 11
0 321 0 0 0 0 0 0 0 0
1
0
0 0 21360 270
2 5V
-6 -21 8 -13
3 V60
-9 -31 12 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
5866 0 0
2
5.89983e-315 5.44228e-315
0
13 Logic Switch~
5 2714 1680 0 10 11
0 320 0 0 0 0 0 0 0 0
1
0
0 0 21360 270
2 5V
-6 -21 8 -13
3 V59
-9 -31 12 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3541 0 0
2
5.89983e-315 5.44487e-315
0
13 Logic Switch~
5 2679 1680 0 10 11
0 319 0 0 0 0 0 0 0 0
1
0
0 0 21360 270
2 5V
-6 -21 8 -13
3 V58
-9 -31 12 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
8710 0 0
2
5.89983e-315 5.44746e-315
0
13 Logic Switch~
5 2392 1688 0 1 11
0 327
0
0 0 21360 270
2 0V
-6 -21 8 -13
3 V57
-9 -31 12 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
8575 0 0
2
5.89983e-315 5.45005e-315
0
13 Logic Switch~
5 2427 1688 0 1 11
0 328
0
0 0 21360 270
2 0V
-6 -21 8 -13
3 V56
-9 -31 12 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
6774 0 0
2
5.89983e-315 5.45264e-315
0
13 Logic Switch~
5 2458 1688 0 1 11
0 329
0
0 0 21360 270
2 0V
-6 -21 8 -13
3 V55
-9 -31 12 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
4257 0 0
2
5.89983e-315 5.45523e-315
0
13 Logic Switch~
5 2491 1688 0 1 11
0 330
0
0 0 21360 270
2 0V
-6 -21 8 -13
3 V54
-9 -31 12 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
5226 0 0
2
5.89983e-315 5.45782e-315
0
13 Logic Switch~
5 2775 1996 0 10 11
0 306 0 0 0 0 0 0 0 0
1
0
0 0 21360 270
2 5V
-6 -21 8 -13
3 V53
-9 -31 12 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
4273 0 0
2
5.89983e-315 5.46041e-315
0
13 Logic Switch~
5 2742 1996 0 10 11
0 305 0 0 0 0 0 0 0 0
1
0
0 0 21360 270
2 5V
-6 -21 8 -13
3 V52
-9 -31 12 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
7945 0 0
2
5.89983e-315 5.463e-315
0
13 Logic Switch~
5 2711 1996 0 1 11
0 304
0
0 0 21360 270
2 0V
-6 -21 8 -13
3 V51
-9 -31 12 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
523 0 0
2
5.89983e-315 5.46559e-315
0
13 Logic Switch~
5 2676 1996 0 1 11
0 303
0
0 0 21360 270
2 0V
-6 -21 8 -13
3 V50
-9 -31 12 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
7617 0 0
2
5.89983e-315 5.46818e-315
0
13 Logic Switch~
5 2389 2004 0 10 11
0 311 0 0 0 0 0 0 0 0
1
0
0 0 21360 270
2 5V
-6 -21 8 -13
3 V49
-9 -31 12 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3526 0 0
2
5.89983e-315 5.47077e-315
0
13 Logic Switch~
5 2424 2004 0 1 11
0 312
0
0 0 21360 270
2 0V
-6 -21 8 -13
3 V48
-9 -31 12 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
3556 0 0
2
5.89983e-315 5.47207e-315
0
13 Logic Switch~
5 2455 2004 0 1 11
0 313
0
0 0 21360 270
2 0V
-6 -21 8 -13
3 V47
-9 -31 12 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
9943 0 0
2
5.89983e-315 5.47336e-315
0
13 Logic Switch~
5 2488 2004 0 10 11
0 314 0 0 0 0 0 0 0 0
1
0
0 0 21360 270
2 5V
-6 -21 8 -13
3 V46
-9 -31 12 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
8750 0 0
2
5.89983e-315 5.47466e-315
0
13 Logic Switch~
5 2776 2332 0 10 11
0 290 0 0 0 0 0 0 0 0
1
0
0 0 21360 270
2 5V
-6 -21 8 -13
3 V45
-9 -31 12 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3208 0 0
2
5.89983e-315 5.47595e-315
0
13 Logic Switch~
5 2743 2332 0 1 11
0 289
0
0 0 21360 270
2 0V
-6 -21 8 -13
3 V44
-9 -31 12 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
6594 0 0
2
5.89983e-315 5.47725e-315
0
13 Logic Switch~
5 2712 2332 0 1 11
0 288
0
0 0 21360 270
2 0V
-6 -21 8 -13
3 V43
-9 -31 12 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
324 0 0
2
5.89983e-315 5.47854e-315
0
13 Logic Switch~
5 2677 2332 0 10 11
0 287 0 0 0 0 0 0 0 0
1
0
0 0 21360 270
2 5V
-6 -21 8 -13
3 V42
-9 -31 12 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
7980 0 0
2
5.89983e-315 5.47984e-315
0
13 Logic Switch~
5 2390 2340 0 10 11
0 295 0 0 0 0 0 0 0 0
1
0
0 0 21360 270
2 5V
-6 -21 8 -13
3 V41
-9 -31 12 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
5129 0 0
2
5.89983e-315 5.48113e-315
0
13 Logic Switch~
5 2425 2340 0 10 11
0 296 0 0 0 0 0 0 0 0
1
0
0 0 21360 270
2 5V
-6 -21 8 -13
3 V40
-9 -31 12 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
6641 0 0
2
5.89983e-315 5.48243e-315
0
13 Logic Switch~
5 2456 2340 0 10 11
0 297 0 0 0 0 0 0 0 0
1
0
0 0 21360 270
2 5V
-6 -21 8 -13
3 V39
-9 -31 12 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
8473 0 0
2
5.89983e-315 5.48372e-315
0
13 Logic Switch~
5 2489 2340 0 1 11
0 298
0
0 0 21360 270
2 0V
-6 -21 8 -13
3 V38
-9 -31 12 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
3989 0 0
2
5.89983e-315 5.48502e-315
0
13 Logic Switch~
5 2481 1066 0 1 11
0 346
0
0 0 21360 270
2 0V
-6 -21 8 -13
3 V37
-9 -31 12 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
3603 0 0
2
5.89983e-315 5.48631e-315
0
13 Logic Switch~
5 2448 1066 0 1 11
0 345
0
0 0 21360 270
2 0V
-6 -21 8 -13
3 V36
-9 -31 12 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
9162 0 0
2
5.89983e-315 5.48761e-315
0
13 Logic Switch~
5 2417 1066 0 10 11
0 344 0 0 0 0 0 0 0 0
1
0
0 0 21360 270
2 5V
-6 -21 8 -13
3 V35
-9 -31 12 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
8123 0 0
2
5.89983e-315 5.4889e-315
0
13 Logic Switch~
5 2382 1066 0 10 11
0 343 0 0 0 0 0 0 0 0
1
0
0 0 21360 270
2 5V
-6 -21 8 -13
3 V34
-9 -31 12 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
4518 0 0
2
5.89983e-315 5.4902e-315
0
13 Logic Switch~
5 2669 1058 0 10 11
0 335 0 0 0 0 0 0 0 0
1
0
0 0 21360 270
2 5V
-6 -21 8 -13
3 V33
-9 -31 12 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3901 0 0
2
5.89983e-315 5.49149e-315
0
13 Logic Switch~
5 2704 1058 0 10 11
0 336 0 0 0 0 0 0 0 0
1
0
0 0 21360 270
2 5V
-6 -21 8 -13
3 V32
-9 -31 12 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
8682 0 0
2
5.89983e-315 5.49279e-315
0
13 Logic Switch~
5 2735 1058 0 10 11
0 337 0 0 0 0 0 0 0 0
1
0
0 0 21360 270
2 5V
-6 -21 8 -13
3 V31
-9 -31 12 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
9523 0 0
2
5.89983e-315 5.49408e-315
0
13 Logic Switch~
5 2768 1058 0 10 11
0 338 0 0 0 0 0 0 0 0
1
0
0 0 21360 270
2 5V
-6 -21 8 -13
3 V30
-9 -31 12 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
5998 0 0
2
5.89983e-315 5.49538e-315
0
13 Logic Switch~
5 2480 730 0 1 11
0 358
0
0 0 21360 270
2 0V
-6 -21 8 -13
3 V29
-9 -31 12 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
4812 0 0
2
5.89983e-315 5.49667e-315
0
13 Logic Switch~
5 2447 730 0 10 11
0 357 0 0 0 0 0 0 0 0
1
0
0 0 21360 270
2 5V
-6 -21 8 -13
3 V28
-9 -31 12 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
7277 0 0
2
5.89983e-315 5.49797e-315
0
13 Logic Switch~
5 2416 730 0 1 11
0 356
0
0 0 21360 270
2 0V
-6 -21 8 -13
3 V27
-9 -31 12 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3564 0 0
2
5.89983e-315 5.49926e-315
0
13 Logic Switch~
5 2381 730 0 10 11
0 355 0 0 0 0 0 0 0 0
1
0
0 0 21360 270
2 5V
-6 -21 8 -13
3 V26
-9 -31 12 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
9696 0 0
2
5.89983e-315 5.50056e-315
0
13 Logic Switch~
5 2668 722 0 1 11
0 347
0
0 0 21360 270
2 0V
-6 -21 8 -13
3 V25
-9 -31 12 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
6303 0 0
2
5.89983e-315 5.50185e-315
0
13 Logic Switch~
5 2703 722 0 1 11
0 348
0
0 0 21360 270
2 0V
-6 -21 8 -13
3 V24
-9 -31 12 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
6155 0 0
2
5.89983e-315 5.50315e-315
0
13 Logic Switch~
5 2734 722 0 1 11
0 349
0
0 0 21360 270
2 0V
-6 -21 8 -13
3 V23
-9 -31 12 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
3180 0 0
2
5.89983e-315 5.50444e-315
0
13 Logic Switch~
5 2767 722 0 1 11
0 350
0
0 0 21360 270
2 0V
-6 -21 8 -13
3 V22
-9 -31 12 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
7733 0 0
2
5.89983e-315 5.50574e-315
0
13 Logic Switch~
5 2760 139 0 10 11
0 366 0 0 0 0 0 0 0 0
1
0
0 0 21360 270
2 5V
-6 -21 8 -13
3 V13
-9 -31 12 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
674 0 0
2
5.89983e-315 5.50703e-315
0
13 Logic Switch~
5 2727 139 0 1 11
0 365
0
0 0 21360 270
2 0V
-6 -21 8 -13
3 V12
-9 -31 12 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
3341 0 0
2
5.89983e-315 5.50833e-315
0
13 Logic Switch~
5 2696 139 0 1 11
0 364
0
0 0 21360 270
2 0V
-6 -21 8 -13
3 V11
-9 -31 12 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
7159 0 0
2
5.89983e-315 5.50963e-315
0
13 Logic Switch~
5 2661 139 0 10 11
0 363 0 0 0 0 0 0 0 0
1
0
0 0 21360 270
2 5V
-6 -21 8 -13
3 V10
-9 -31 12 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3833 0 0
2
5.89983e-315 5.51092e-315
0
13 Logic Switch~
5 2374 147 0 1 11
0 371
0
0 0 21360 270
2 0V
-6 -21 8 -13
2 V6
-6 -31 8 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
4828 0 0
2
5.89983e-315 5.51222e-315
0
13 Logic Switch~
5 2409 147 0 10 11
0 372 0 0 0 0 0 0 0 0
1
0
0 0 21360 270
2 5V
-6 -21 8 -13
2 V7
-6 -31 8 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3263 0 0
2
5.89983e-315 5.51286e-315
0
13 Logic Switch~
5 2440 147 0 1 11
0 373
0
0 0 21360 270
2 0V
-6 -21 8 -13
2 V8
-6 -31 8 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
3250 0 0
2
5.89983e-315 5.51351e-315
0
13 Logic Switch~
5 2473 147 0 10 11
0 374 0 0 0 0 0 0 0 0
1
0
0 0 21360 270
2 5V
-6 -21 8 -13
2 V9
-6 -31 8 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3550 0 0
2
5.89983e-315 5.51416e-315
0
13 Logic Switch~
5 135 369 0 10 11
0 384 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-5 -16 9 -8
2 V1
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
9418 0 0
2
44331.3 0
0
13 Logic Switch~
5 135 486 0 1 11
0 391
0
0 0 21360 0
2 0V
-5 -16 9 -8
2 V1
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
335 0 0
2
44331.3 1
0
13 Logic Switch~
5 135 538 0 10 11
0 390 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V2
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
9178 0 0
2
44331.3 2
0
13 Logic Switch~
5 136 584 0 1 11
0 389
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V3
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
4802 0 0
2
44331.3 3
0
13 Logic Switch~
5 136 631 0 10 11
0 388 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V4
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
4114 0 0
2
44331.3 4
0
9 Inverter~
13 2848 2547 0 2 22
0 4 106
0
0 0 624 512
6 74LS04
-21 -19 21 -11
4 U95E
-8 -20 20 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 11 10 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 5 36 0
1 U
3439 0 0
2
5.89983e-315 5.51481e-315
0
9 Inverter~
13 2845 2220 0 2 22
0 5 107
0
0 0 624 512
6 74LS04
-21 -19 21 -11
4 U95D
-8 -20 20 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 9 8 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 4 36 0
1 U
8948 0 0
2
5.89983e-315 5.51545e-315
0
9 Inverter~
13 2844 1899 0 2 22
0 6 109
0
0 0 624 512
6 74LS04
-21 -19 21 -11
4 U95C
-8 -20 20 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 5 6 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 3 36 0
1 U
4509 0 0
2
5.89983e-315 5.5161e-315
0
9 Inverter~
13 2853 1594 0 2 22
0 7 110
0
0 0 624 512
6 74LS04
-21 -19 21 -11
4 U95B
-8 -20 20 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 3 4 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 2 36 0
1 U
5161 0 0
2
5.89983e-315 5.51675e-315
0
14 Logic Display~
6 1708 1575 0 1 2
10 12
0
0 0 53856 0
6 100MEG
3 -16 45 -8
4 L147
-13 -21 15 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
8614 0 0
2
5.89983e-315 5.5174e-315
0
14 Logic Display~
6 1724 1575 0 1 2
10 11
0
0 0 53856 0
6 100MEG
3 -16 45 -8
4 L146
-13 -21 15 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
661 0 0
2
5.89983e-315 5.51804e-315
0
14 Logic Display~
6 1740 1575 0 1 2
10 10
0
0 0 53856 0
6 100MEG
3 -16 45 -8
4 L145
-13 -21 15 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
8325 0 0
2
5.89983e-315 5.51869e-315
0
14 Logic Display~
6 1756 1575 0 1 2
10 9
0
0 0 53856 0
6 100MEG
3 -16 45 -8
4 L144
-13 -21 15 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
335 0 0
2
5.89983e-315 5.51934e-315
0
14 Logic Display~
6 1706 1054 0 1 2
10 16
0
0 0 53856 0
6 100MEG
3 -16 45 -8
4 L143
-13 -21 15 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
4239 0 0
2
5.89983e-315 5.51999e-315
0
14 Logic Display~
6 1722 1054 0 1 2
10 15
0
0 0 53856 0
6 100MEG
3 -16 45 -8
4 L142
-13 -21 15 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
49 0 0
2
5.89983e-315 5.52063e-315
0
14 Logic Display~
6 1738 1054 0 1 2
10 14
0
0 0 53856 0
6 100MEG
3 -16 45 -8
4 L141
-13 -21 15 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
9471 0 0
2
5.89983e-315 5.52128e-315
0
14 Logic Display~
6 1754 1054 0 1 2
10 13
0
0 0 53856 0
6 100MEG
3 -16 45 -8
4 L140
-13 -21 15 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3808 0 0
2
5.89983e-315 5.52193e-315
0
14 Logic Display~
6 1701 662 0 1 2
10 20
0
0 0 53856 0
6 100MEG
3 -16 45 -8
4 L139
-13 -21 15 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
9213 0 0
2
5.89983e-315 5.52258e-315
0
14 Logic Display~
6 1717 662 0 1 2
10 19
0
0 0 53856 0
6 100MEG
3 -16 45 -8
4 L138
-13 -21 15 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3504 0 0
2
5.89983e-315 5.52322e-315
0
14 Logic Display~
6 1733 662 0 1 2
10 18
0
0 0 53856 0
6 100MEG
3 -16 45 -8
4 L137
-13 -21 15 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
4873 0 0
2
5.89983e-315 5.52387e-315
0
14 Logic Display~
6 1749 662 0 1 2
10 17
0
0 0 53856 0
6 100MEG
3 -16 45 -8
3 L92
-9 -21 12 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
65 0 0
2
5.89983e-315 5.52452e-315
0
14 Logic Display~
6 1743 255 0 1 2
10 21
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L1
-6 -21 8 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3246 0 0
2
5.89983e-315 5.52517e-315
0
14 Logic Display~
6 1727 255 0 1 2
10 22
0
0 0 53856 0
6 100MEG
3 -16 45 -8
3 L89
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
5176 0 0
2
5.89983e-315 5.52581e-315
0
14 Logic Display~
6 1711 255 0 1 2
10 23
0
0 0 53856 0
6 100MEG
3 -16 45 -8
3 L90
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3796 0 0
2
5.89983e-315 5.52646e-315
0
14 Logic Display~
6 1695 255 0 1 2
10 24
0
0 0 53856 0
6 100MEG
3 -16 45 -8
3 L91
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3359 0 0
2
5.89983e-315 5.52711e-315
0
14 Logic Display~
6 1277 1580 0 1 2
10 28
0
0 0 53856 0
6 100MEG
3 -16 45 -8
4 L136
-13 -21 15 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
8339 0 0
2
5.89983e-315 5.52776e-315
0
14 Logic Display~
6 1293 1580 0 1 2
10 27
0
0 0 53856 0
6 100MEG
3 -16 45 -8
4 L135
-13 -21 15 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3578 0 0
2
5.89983e-315 5.52841e-315
0
14 Logic Display~
6 1309 1580 0 1 2
10 26
0
0 0 53856 0
6 100MEG
3 -16 45 -8
4 L134
-13 -21 15 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
4575 0 0
2
5.89983e-315 5.52905e-315
0
14 Logic Display~
6 1325 1580 0 1 2
10 25
0
0 0 53856 0
6 100MEG
3 -16 45 -8
4 L133
-13 -21 15 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
6878 0 0
2
5.89983e-315 5.5297e-315
0
14 Logic Display~
6 1270 1060 0 1 2
10 32
0
0 0 53856 0
6 100MEG
3 -16 45 -8
4 L132
-13 -21 15 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
8570 0 0
2
5.89983e-315 5.53035e-315
0
14 Logic Display~
6 1286 1060 0 1 2
10 31
0
0 0 53856 0
6 100MEG
3 -16 45 -8
4 L131
-13 -21 15 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3708 0 0
2
5.89983e-315 5.531e-315
0
14 Logic Display~
6 1302 1060 0 1 2
10 30
0
0 0 53856 0
6 100MEG
3 -16 45 -8
4 L130
-13 -21 15 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3251 0 0
2
5.89983e-315 5.53164e-315
0
14 Logic Display~
6 1318 1060 0 1 2
10 29
0
0 0 53856 0
6 100MEG
3 -16 45 -8
4 L129
-13 -21 15 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3597 0 0
2
5.89983e-315 5.53229e-315
0
14 Logic Display~
6 1261 667 0 1 2
10 36
0
0 0 53856 0
6 100MEG
3 -16 45 -8
4 L128
-13 -21 15 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
4380 0 0
2
5.89983e-315 5.53294e-315
0
14 Logic Display~
6 1277 667 0 1 2
10 35
0
0 0 53856 0
6 100MEG
3 -16 45 -8
4 L127
-13 -21 15 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
4808 0 0
2
5.89983e-315 5.53359e-315
0
14 Logic Display~
6 1293 667 0 1 2
10 34
0
0 0 53856 0
6 100MEG
3 -16 45 -8
4 L126
-13 -21 15 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
7106 0 0
2
5.89983e-315 5.53423e-315
0
14 Logic Display~
6 1309 667 0 1 2
10 33
0
0 0 53856 0
6 100MEG
3 -16 45 -8
4 L125
-13 -21 15 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
345 0 0
2
5.89983e-315 5.53488e-315
0
14 Logic Display~
6 1305 256 0 1 2
10 37
0
0 0 53856 0
6 100MEG
3 -16 45 -8
4 L124
-13 -21 15 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
5150 0 0
2
5.89983e-315 5.53553e-315
0
14 Logic Display~
6 1289 256 0 1 2
10 38
0
0 0 53856 0
6 100MEG
3 -16 45 -8
4 L123
-13 -21 15 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
5481 0 0
2
5.89983e-315 5.53618e-315
0
14 Logic Display~
6 1273 256 0 1 2
10 39
0
0 0 53856 0
6 100MEG
3 -16 45 -8
4 L122
-13 -21 15 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
6899 0 0
2
5.89983e-315 5.53682e-315
0
14 Logic Display~
6 1257 256 0 1 2
10 40
0
0 0 53856 0
6 100MEG
3 -16 45 -8
4 L121
-13 -21 15 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
6995 0 0
2
5.89983e-315 5.53747e-315
0
8 2-In OR~
219 1646 1753 0 3 22
0 42 43 115
0
0 0 624 90
6 74LS32
-21 -24 21 -16
4 U96A
-12 -5 16 3
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 37 0
1 U
3497 0 0
2
5.89983e-315 5.53812e-315
0
8 2-In OR~
219 1648 1221 0 3 22
0 46 45 44
0
0 0 624 90
6 74LS32
-21 -24 21 -16
4 U93D
-12 -5 16 3
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 34 0
1 U
4890 0 0
2
5.89983e-315 5.53877e-315
0
8 2-In OR~
219 1642 802 0 3 22
0 49 48 116
0
0 0 624 90
6 74LS32
-21 -24 21 -16
4 U93C
-12 -5 16 3
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 9 10 8 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 34 0
1 U
4995 0 0
2
5.89983e-315 5.53941e-315
0
9 Inverter~
13 1502 1936 0 2 22
0 406 407
0
0 0 624 0
6 74LS04
-21 -19 21 -11
4 U95A
-14 -20 14 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 512 6 1 36 0
1 U
3337 0 0
2
5.89983e-315 5.54006e-315
0
8 2-In OR~
219 1646 389 0 3 22
0 59 58 47
0
0 0 624 90
6 74LS32
-21 -24 21 -16
4 U93B
-12 -5 16 3
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 34 0
1 U
548 0 0
2
5.89983e-315 5.54071e-315
0
14 Logic Display~
6 948 676 0 1 2
10 61
0
0 0 53856 0
6 100MEG
3 -16 45 -8
3 L76
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
5680 0 0
2
5.89983e-315 5.54136e-315
0
14 Logic Display~
6 939 277 0 1 2
10 62
0
0 0 53856 0
6 100MEG
3 -16 45 -8
3 L73
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3208 0 0
2
5.89983e-315 5.542e-315
0
14 Logic Display~
6 1583 1744 0 1 2
10 64
0
0 0 53856 180
6 100MEG
3 -16 45 -8
4 L120
-5 18 23 26
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
4420 0 0
2
5.89983e-315 5.54265e-315
0
14 Logic Display~
6 1599 1744 0 1 2
10 63
0
0 0 53856 180
6 100MEG
3 -16 45 -8
4 L119
8 0 36 8
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
5529 0 0
2
5.89983e-315 5.5433e-315
0
14 Logic Display~
6 1567 1744 0 1 2
10 65
0
0 0 53856 180
6 100MEG
3 -16 45 -8
4 L118
-13 18 15 26
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
8579 0 0
2
5.89983e-315 5.54395e-315
0
14 Logic Display~
6 1551 1744 0 1 2
10 66
0
0 0 53856 180
6 100MEG
3 -16 45 -8
4 L117
-22 18 6 26
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
5723 0 0
2
5.89983e-315 5.54459e-315
0
14 Logic Display~
6 1393 1744 0 1 2
10 68
0
0 0 53856 180
6 100MEG
3 -16 45 -8
4 L116
-5 18 23 26
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3325 0 0
2
5.89983e-315 5.54524e-315
0
14 Logic Display~
6 1409 1744 0 1 2
10 67
0
0 0 53856 180
6 100MEG
3 -16 45 -8
4 L115
8 0 36 8
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3552 0 0
2
5.89983e-315 5.54589e-315
0
14 Logic Display~
6 1377 1744 0 1 2
10 69
0
0 0 53856 180
6 100MEG
3 -16 45 -8
4 L114
-13 18 15 26
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
8709 0 0
2
5.89983e-315 5.54654e-315
0
14 Logic Display~
6 1361 1744 0 1 2
10 70
0
0 0 53856 180
6 100MEG
3 -16 45 -8
4 L113
-22 18 6 26
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3346 0 0
2
5.89983e-315 5.54719e-315
0
14 Logic Display~
6 1581 1211 0 1 2
10 72
0
0 0 53856 180
6 100MEG
3 -16 45 -8
4 L112
-5 18 23 26
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3220 0 0
2
5.89983e-315 5.54783e-315
0
14 Logic Display~
6 1597 1211 0 1 2
10 71
0
0 0 53856 180
6 100MEG
3 -16 45 -8
4 L111
8 0 36 8
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
4894 0 0
2
5.89983e-315 5.54848e-315
0
14 Logic Display~
6 1565 1211 0 1 2
10 73
0
0 0 53856 180
6 100MEG
3 -16 45 -8
4 L110
-13 18 15 26
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
8598 0 0
2
5.89983e-315 5.54913e-315
0
14 Logic Display~
6 1549 1211 0 1 2
10 74
0
0 0 53856 180
6 100MEG
3 -16 45 -8
4 L109
-22 18 6 26
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
4222 0 0
2
5.89983e-315 5.54978e-315
0
14 Logic Display~
6 1386 1212 0 1 2
10 76
0
0 0 53856 180
6 100MEG
3 -16 45 -8
4 L108
-5 18 23 26
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
6818 0 0
2
5.89983e-315 5.55042e-315
0
14 Logic Display~
6 1402 1212 0 1 2
10 75
0
0 0 53856 180
6 100MEG
3 -16 45 -8
4 L107
8 0 36 8
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
783 0 0
2
5.89983e-315 5.55107e-315
0
14 Logic Display~
6 1370 1212 0 1 2
10 77
0
0 0 53856 180
6 100MEG
3 -16 45 -8
4 L106
-13 18 15 26
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
7884 0 0
2
5.89983e-315 5.55172e-315
0
14 Logic Display~
6 1354 1212 0 1 2
10 78
0
0 0 53856 180
6 100MEG
3 -16 45 -8
4 L105
-22 18 6 26
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
8282 0 0
2
5.89983e-315 5.55237e-315
0
14 Logic Display~
6 1576 800 0 1 2
10 80
0
0 0 53856 180
6 100MEG
3 -16 45 -8
4 L104
-5 18 23 26
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
6937 0 0
2
5.89983e-315 5.55301e-315
0
14 Logic Display~
6 1592 800 0 1 2
10 79
0
0 0 53856 180
6 100MEG
3 -16 45 -8
4 L103
8 0 36 8
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3682 0 0
2
5.89983e-315 5.55366e-315
0
14 Logic Display~
6 1560 800 0 1 2
10 81
0
0 0 53856 180
6 100MEG
3 -16 45 -8
4 L102
-13 18 15 26
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
8332 0 0
2
5.89983e-315 5.55398e-315
0
14 Logic Display~
6 1544 800 0 1 2
10 82
0
0 0 53856 180
6 100MEG
3 -16 45 -8
4 L101
-22 18 6 26
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3772 0 0
2
5.89983e-315 5.55431e-315
0
14 Logic Display~
6 1570 382 0 1 2
10 84
0
0 0 53856 180
6 100MEG
3 -16 45 -8
4 L100
-5 18 23 26
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
4564 0 0
2
5.89983e-315 5.55463e-315
0
14 Logic Display~
6 1586 382 0 1 2
10 83
0
0 0 53856 180
6 100MEG
3 -16 45 -8
3 L99
11 0 32 8
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
5280 0 0
2
5.89983e-315 5.55496e-315
0
14 Logic Display~
6 1554 382 0 1 2
10 85
0
0 0 53856 180
6 100MEG
3 -16 45 -8
3 L98
-10 18 11 26
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
4934 0 0
2
5.89983e-315 5.55528e-315
0
14 Logic Display~
6 1538 382 0 1 2
10 86
0
0 0 53856 180
6 100MEG
3 -16 45 -8
3 L97
-19 18 2 26
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
390 0 0
2
5.89983e-315 5.5556e-315
0
14 Logic Display~
6 1373 380 0 1 2
10 88
0
0 0 53856 180
6 100MEG
3 -16 45 -8
3 L96
-2 18 19 26
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
45 0 0
2
5.89983e-315 5.55593e-315
0
14 Logic Display~
6 1389 380 0 1 2
10 87
0
0 0 53856 180
6 100MEG
3 -16 45 -8
3 L95
11 0 32 8
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
7163 0 0
2
5.89983e-315 5.55625e-315
0
14 Logic Display~
6 1357 380 0 1 2
10 89
0
0 0 53856 180
6 100MEG
3 -16 45 -8
3 L94
-10 18 11 26
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
4130 0 0
2
5.89983e-315 5.55657e-315
0
14 Logic Display~
6 1341 380 0 1 2
10 90
0
0 0 53856 180
6 100MEG
3 -16 45 -8
3 L93
-19 18 2 26
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
7512 0 0
2
5.89983e-315 5.5569e-315
0
14 Logic Display~
6 1348 802 0 1 2
10 94
0
0 0 53856 180
6 100MEG
3 -16 45 -8
3 L85
-19 18 2 26
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
7351 0 0
2
5.89983e-315 5.55722e-315
0
14 Logic Display~
6 1363 802 0 1 2
10 93
0
0 0 53856 180
6 100MEG
3 -16 45 -8
3 L86
-10 18 11 26
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3114 0 0
2
5.89983e-315 5.55755e-315
0
14 Logic Display~
6 1394 802 0 1 2
10 91
0
0 0 53856 180
6 100MEG
3 -16 45 -8
3 L88
11 0 32 8
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3304 0 0
2
5.89983e-315 5.55787e-315
0
14 Logic Display~
6 1378 802 0 1 2
10 92
0
0 0 53856 180
6 100MEG
3 -16 45 -8
3 L87
-2 18 19 26
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3640 0 0
2
5.89983e-315 5.55819e-315
0
14 Logic Display~
6 1294 1677 0 1 2
10 95
0
0 0 53856 0
6 100MEG
3 -16 45 -8
3 L84
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
739 0 0
2
5.89983e-315 5.55852e-315
0
14 Logic Display~
6 1142 1585 0 1 2
10 96
0
0 0 53856 0
6 100MEG
3 -16 45 -8
3 L83
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
4482 0 0
2
5.89983e-315 5.55884e-315
0
14 Logic Display~
6 986 1588 0 1 2
10 97
0
0 0 53856 0
6 100MEG
3 -16 45 -8
3 L82
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
6605 0 0
2
5.89983e-315 5.55917e-315
0
14 Logic Display~
6 1278 1122 0 1 2
10 98
0
0 0 53856 0
6 100MEG
3 -16 45 -8
3 L81
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
7726 0 0
2
5.89983e-315 5.55949e-315
0
14 Logic Display~
6 967 1050 0 1 2
10 99
0
0 0 53856 0
6 100MEG
3 -16 45 -8
3 L80
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
9904 0 0
2
5.89983e-315 5.55981e-315
0
14 Logic Display~
6 1144 1055 0 1 2
10 100
0
0 0 53856 0
6 100MEG
3 -16 45 -8
3 L79
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
4780 0 0
2
5.89983e-315 5.56014e-315
0
14 Logic Display~
6 1256 740 0 1 2
10 101
0
0 0 53856 0
6 100MEG
3 -16 45 -8
3 L78
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
4251 0 0
2
5.89983e-315 5.56046e-315
0
14 Logic Display~
6 1120 678 0 1 2
10 102
0
0 0 53856 0
6 100MEG
3 -16 45 -8
3 L77
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
6909 0 0
2
5.89983e-315 5.56078e-315
0
14 Logic Display~
6 1257 338 0 1 2
10 103
0
0 0 53856 0
6 100MEG
3 -16 45 -8
3 L75
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3348 0 0
2
5.89983e-315 5.56111e-315
0
14 Logic Display~
6 1111 284 0 1 2
10 104
0
0 0 53856 0
6 100MEG
3 -16 45 -8
3 L74
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
4560 0 0
2
5.89983e-315 5.56143e-315
0
8 2-In OR~
219 1035 1521 0 3 22
0 106 105 111
0
0 0 624 270
6 74LS32
-21 -24 21 -16
4 U93A
-10 -8 18 0
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 34 0
1 U
3137 0 0
2
44331.3 5
0
8 2-In OR~
219 1023 988 0 3 22
0 107 108 112
0
0 0 624 270
6 74LS32
-21 -24 21 -16
4 U89D
-10 -8 18 0
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 30 0
1 U
9152 0 0
2
44331.3 6
0
8 2-In OR~
219 1005 597 0 3 22
0 109 8 113
0
0 0 624 270
6 74LS32
-21 -24 21 -16
4 U89C
-10 -8 18 0
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 9 10 8 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 30 0
1 U
3390 0 0
2
44331.3 7
0
8 2-In OR~
219 1002 202 0 3 22
0 110 60 114
0
0 0 624 270
6 74LS32
-21 -24 21 -16
4 U89B
-10 -8 18 0
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 30 0
1 U
43 0 0
2
44331.3 8
0
10 Buffer 3S~
219 1023 1629 0 3 22
0 117 115 118
0
0 0 624 0
8 BUFFER3S
-27 -51 29 -43
4 U92B
-11 -12 17 -4
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
0
22

0 5 4 6 2 1 3 5 4 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 33 0
1 U
3347 0 0
2
44331.3 9
0
10 Buffer 3S~
219 1037 1584 0 3 22
0 111 115 119
0
0 0 624 0
8 BUFFER3S
-27 -51 29 -43
4 U92A
-14 -20 14 -12
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
0
22

0 2 1 3 2 1 3 5 4 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 33 0
1 U
8673 0 0
2
44331.3 10
0
10 Buffer 3S~
219 1023 1099 0 3 22
0 117 44 120
0
0 0 624 0
8 BUFFER3S
-27 -51 29 -43
4 U91D
-11 -12 17 -4
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
0
22

0 12 13 11 2 1 3 5 4 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 32 0
1 U
3232 0 0
2
44331.3 11
0
10 Buffer 3S~
219 1037 1054 0 3 22
0 112 44 121
0
0 0 624 0
8 BUFFER3S
-27 -51 29 -43
4 U91C
-14 -20 14 -12
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
0
22

0 9 10 8 2 1 3 5 4 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 32 0
1 U
8598 0 0
2
44331.3 12
0
10 Buffer 3S~
219 999 722 0 3 22
0 117 116 122
0
0 0 624 0
8 BUFFER3S
-27 -51 29 -43
4 U91B
-11 -12 17 -4
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
0
22

0 5 4 6 2 1 3 5 4 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 32 0
1 U
8765 0 0
2
44331.3 13
0
10 Buffer 3S~
219 1013 677 0 3 22
0 113 116 123
0
0 0 624 0
8 BUFFER3S
-27 -51 29 -43
4 U91A
-14 -20 14 -12
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
0
22

0 2 1 3 2 1 3 5 4 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 32 0
1 U
4481 0 0
2
44331.3 14
0
10 Buffer 3S~
219 1003 283 0 3 22
0 114 47 125
0
0 0 624 0
8 BUFFER3S
-27 -51 29 -43
4 U90B
-14 -20 14 -12
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
0
22

0 5 4 6 2 1 3 5 4 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 31 0
1 U
7314 0 0
2
44331.3 15
0
10 Buffer 3S~
219 989 328 0 3 22
0 117 47 124
0
0 0 624 0
8 BUFFER3S
-27 -51 29 -43
4 U90A
-11 -12 17 -4
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
0
22

0 2 1 3 2 1 3 5 4 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 31 0
1 U
3331 0 0
2
44331.3 16
0
10 Buffer 3S~
219 877 1632 0 3 22
0 117 115 127
0
0 0 624 0
8 BUFFER3S
-27 -51 29 -43
4 U88A
-11 -12 17 -4
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
0
22

0 2 1 3 2 1 3 5 4 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 29 0
1 U
3179 0 0
2
5.89983e-315 5.56176e-315
0
10 Buffer 3S~
219 877 1587 0 3 22
0 126 115 128
0
0 0 624 0
8 BUFFER3S
-27 -51 29 -43
4 U87D
-14 -20 14 -12
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
0
22

0 12 13 11 2 1 3 5 4 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 28 0
1 U
7409 0 0
2
5.89983e-315 5.56208e-315
0
10 Buffer 3S~
219 865 1096 0 3 22
0 117 44 130
0
0 0 624 0
8 BUFFER3S
-27 -51 29 -43
4 U87C
-11 -12 17 -4
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
0
22

0 9 10 8 2 1 3 5 4 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 28 0
1 U
3276 0 0
2
5.89983e-315 5.5624e-315
0
10 Buffer 3S~
219 865 1051 0 3 22
0 129 44 131
0
0 0 624 0
8 BUFFER3S
-27 -51 29 -43
4 U87B
-14 -20 14 -12
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
0
22

0 5 4 6 2 1 3 5 4 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 28 0
1 U
3169 0 0
2
5.89983e-315 5.56273e-315
0
10 Buffer 3S~
219 843 719 0 3 22
0 117 116 133
0
0 0 624 0
8 BUFFER3S
-27 -51 29 -43
4 U87A
-11 -12 17 -4
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
0
22

0 2 1 3 2 1 3 5 4 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 28 0
1 U
3896 0 0
2
5.89983e-315 5.56305e-315
0
10 Buffer 3S~
219 843 674 0 3 22
0 132 116 134
0
0 0 624 0
8 BUFFER3S
-27 -51 29 -43
4 U83D
-14 -20 14 -12
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
0
22

0 12 13 11 2 1 3 5 4 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 24 0
1 U
4652 0 0
2
5.89983e-315 5.56337e-315
0
10 Buffer 3S~
219 829 276 0 3 22
0 135 47 137
0
0 0 624 0
8 BUFFER3S
-27 -51 29 -43
4 U83B
-14 -20 14 -12
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
0
22

0 5 4 6 2 1 3 5 4 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 24 0
1 U
3818 0 0
2
5.89983e-315 5.5637e-315
0
10 Buffer 3S~
219 829 321 0 3 22
0 117 47 136
0
0 0 624 0
8 BUFFER3S
-27 -51 29 -43
4 U83C
-11 -12 17 -4
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
0
22

0 9 10 8 2 1 3 5 4 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 24 0
1 U
3839 0 0
2
5.89983e-315 5.56402e-315
0
8 2-In OR~
219 1714 1789 0 3 22
0 139 147 43
0
0 0 624 180
6 74LS32
-21 -24 21 -16
4 U85D
-15 -6 13 2
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 26 0
1 U
5247 0 0
2
44331.3 17
0
8 2-In OR~
219 1714 1827 0 3 22
0 138 146 42
0
0 0 624 180
6 74LS32
-21 -24 21 -16
4 U85C
-19 -7 9 1
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 9 10 8 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 26 0
1 U
7397 0 0
2
44331.3 18
0
8 2-In OR~
219 1746 1296 0 3 22
0 140 150 45
0
0 0 624 180
6 74LS32
-21 -24 21 -16
4 U85A
-19 -7 9 1
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 26 0
1 U
4655 0 0
2
44331.3 19
0
8 2-In OR~
219 1745 1262 0 3 22
0 141 151 46
0
0 0 624 180
6 74LS32
-21 -24 21 -16
4 U85B
-15 -6 13 2
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 26 0
1 U
3124 0 0
2
44331.3 20
0
8 2-In OR~
219 1733 868 0 3 22
0 142 152 48
0
0 0 624 180
6 74LS32
-21 -24 21 -16
4 U84C
-19 -7 9 1
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 9 10 8 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 25 0
1 U
7799 0 0
2
44331.3 21
0
8 2-In OR~
219 1733 833 0 3 22
0 143 153 49
0
0 0 624 180
6 74LS32
-21 -24 21 -16
4 U84D
-15 -6 13 2
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 25 0
1 U
3160 0 0
2
44331.3 22
0
8 2-In OR~
219 1739 453 0 3 22
0 144 154 58
0
0 0 624 180
6 74LS32
-21 -24 21 -16
4 U84B
-19 -7 9 1
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 25 0
1 U
5785 0 0
2
44331.3 23
0
8 2-In OR~
219 1739 418 0 3 22
0 145 155 59
0
0 0 624 180
6 74LS32
-21 -24 21 -16
4 U84A
-15 -6 13 2
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 25 0
1 U
7832 0 0
2
44331.3 24
0
10 Buffer 3S~
219 1643 1574 0 3 22
0 117 115 148
0
0 0 624 512
8 BUFFER3S
-27 -51 29 -43
4 U83A
-14 -20 14 -12
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
0
22

0 2 1 3 2 1 3 5 4 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 24 0
1 U
9266 0 0
2
44331.3 25
0
10 Buffer 3S~
219 1455 1570 0 3 22
0 117 115 149
0
0 0 624 512
8 BUFFER3S
-27 -51 29 -43
4 U81D
-14 -20 14 -12
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
0
22

0 12 13 11 2 1 3 5 4 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 22 0
1 U
4817 0 0
2
44331.3 26
0
10 Buffer 3S~
219 1641 1056 0 3 22
0 117 44 156
0
0 0 624 512
8 BUFFER3S
-27 -51 29 -43
4 U81C
-14 -20 14 -12
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
0
22

0 9 10 8 2 1 3 5 4 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 22 0
1 U
3836 0 0
2
44331.3 27
0
10 Buffer 3S~
219 1444 1054 0 3 22
0 117 44 157
0
0 0 624 512
8 BUFFER3S
-27 -51 29 -43
4 U81B
-14 -20 14 -12
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
0
22

0 5 4 6 2 1 3 5 4 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 22 0
1 U
3293 0 0
2
44331.3 28
0
10 Buffer 3S~
219 1645 661 0 3 22
0 117 116 158
0
0 0 624 512
8 BUFFER3S
-27 -51 29 -43
4 U81A
-14 -20 14 -12
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
0
22

0 2 1 3 2 1 3 5 4 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 22 0
1 U
5310 0 0
2
44331.3 29
0
10 Buffer 3S~
219 1432 662 0 3 22
0 117 116 159
0
0 0 624 512
8 BUFFER3S
-27 -51 29 -43
3 U4D
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
0
22

0 12 13 11 2 1 3 5 4 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 2 0
1 U
3347 0 0
2
44331.3 30
0
10 Buffer 3S~
219 1627 256 0 3 22
0 117 47 160
0
0 0 624 512
8 BUFFER3S
-27 -51 29 -43
3 U4C
-8 -12 13 -4
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
0
22

0 9 10 8 2 1 3 5 4 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 2 0
1 U
4338 0 0
2
44331.3 31
0
10 Buffer 3S~
219 1429 251 0 3 22
0 117 47 161
0
0 0 624 512
8 BUFFER3S
-27 -51 29 -43
3 U4A
-8 -12 13 -4
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
0
22

0 2 1 3 2 1 3 5 4 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 2 0
1 U
5936 0 0
2
44331.3 32
0
5 4001~
219 2921 2496 0 3 22
0 138 139 4
0
0 0 624 180
4 4001
-14 -24 14 -16
4 U79D
-9 -8 19 0
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 9 0
65 0 0 0 4 4 20 0
1 U
6862 0 0
2
5.89983e-315 5.56435e-315
0
5 4001~
219 2921 2166 0 3 22
0 140 141 5
0
0 0 624 180
4 4001
-14 -24 14 -16
4 U79C
-9 -8 19 0
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 8 9 10 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 9 0
65 0 0 0 4 3 20 0
1 U
7453 0 0
2
5.89983e-315 5.56467e-315
0
5 4001~
219 2919 1849 0 3 22
0 142 143 6
0
0 0 624 180
4 4001
-14 -24 14 -16
4 U79B
-9 -8 19 0
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 5 6 4 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 9 0
65 0 0 0 4 2 20 0
1 U
8671 0 0
2
5.89983e-315 5.56499e-315
0
5 4001~
219 2918 1543 0 3 22
0 144 145 7
0
0 0 624 180
4 4001
-14 -24 14 -16
4 U79A
-9 -8 19 0
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 9 0
65 0 0 0 4 1 20 0
1 U
8380 0 0
2
5.89983e-315 5.56532e-315
0
5 4001~
219 2892 1226 0 3 22
0 146 147 105
0
0 0 624 180
4 4001
-14 -24 14 -16
4 U78D
-9 -8 19 0
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 9 0
65 0 0 0 4 4 19 0
1 U
5924 0 0
2
5.89983e-315 5.56564e-315
0
5 4001~
219 2913 889 0 3 22
0 150 151 108
0
0 0 624 180
4 4001
-14 -24 14 -16
4 U78C
-12 -12 16 -4
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 8 9 10 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 9 0
65 0 0 0 4 3 19 0
1 U
8710 0 0
2
5.89983e-315 5.56596e-315
0
5 4001~
219 2904 582 0 3 22
0 152 153 8
0
0 0 624 180
4 4001
-14 -24 14 -16
4 U78B
-9 -8 19 0
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 5 6 4 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 9 0
65 0 0 0 4 2 19 0
1 U
3736 0 0
2
5.89983e-315 5.56629e-315
0
5 4001~
219 2906 295 0 3 22
0 154 155 60
0
0 0 624 180
4 4001
-14 -24 14 -16
4 U78A
-9 -8 19 0
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 9 0
65 0 0 0 4 1 19 0
1 U
710 0 0
2
5.89983e-315 5.56661e-315
0
8 2-In OR~
219 1521 1500 0 3 22
0 166 198 234
0
0 0 624 270
6 74LS32
-21 -24 21 -16
4 U77D
-10 -8 18 0
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 18 0
1 U
4481 0 0
2
5.89983e-315 5.56694e-315
0
8 2-In OR~
219 1620 1501 0 3 22
0 163 195 232
0
0 0 624 270
6 74LS32
-21 -24 21 -16
4 U77C
-10 -8 18 0
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 9 10 8 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 18 0
1 U
4389 0 0
2
5.89983e-315 5.56726e-315
0
8 2-In OR~
219 1587 1501 0 3 22
0 164 196 231
0
0 0 624 270
6 74LS32
-21 -24 21 -16
4 U77B
-10 -8 18 0
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 18 0
1 U
7904 0 0
2
5.89983e-315 5.56758e-315
0
8 2-In OR~
219 1554 1500 0 3 22
0 165 197 233
0
0 0 624 270
6 74LS32
-21 -24 21 -16
4 U77A
-10 -8 18 0
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 18 0
1 U
6267 0 0
2
5.89983e-315 5.56791e-315
0
8 2-In OR~
219 1331 1497 0 3 22
0 170 202 238
0
0 0 624 270
6 74LS32
-21 -24 21 -16
4 U76D
-10 -8 18 0
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 17 0
1 U
3906 0 0
2
5.89983e-315 5.56823e-315
0
8 2-In OR~
219 1430 1498 0 3 22
0 167 199 236
0
0 0 624 270
6 74LS32
-21 -24 21 -16
4 U76C
-10 -8 18 0
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 9 10 8 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 17 0
1 U
4196 0 0
2
5.89983e-315 5.56856e-315
0
8 2-In OR~
219 1397 1498 0 3 22
0 168 200 235
0
0 0 624 270
6 74LS32
-21 -24 21 -16
4 U76B
-10 -8 18 0
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 17 0
1 U
3280 0 0
2
5.89983e-315 5.56888e-315
0
8 2-In OR~
219 1364 1497 0 3 22
0 169 201 237
0
0 0 624 270
6 74LS32
-21 -24 21 -16
4 U76A
-10 -8 18 0
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 17 0
1 U
9832 0 0
2
5.89983e-315 5.5692e-315
0
8 2-In OR~
219 1519 983 0 3 22
0 174 210 242
0
0 0 624 270
6 74LS32
-21 -24 21 -16
4 U75D
-10 -8 18 0
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 16 0
1 U
8677 0 0
2
5.89983e-315 5.56953e-315
0
8 2-In OR~
219 1618 984 0 3 22
0 171 207 240
0
0 0 624 270
6 74LS32
-21 -24 21 -16
4 U75C
-10 -8 18 0
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 9 10 8 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 16 0
1 U
3309 0 0
2
5.89983e-315 5.56985e-315
0
8 2-In OR~
219 1585 984 0 3 22
0 172 208 239
0
0 0 624 270
6 74LS32
-21 -24 21 -16
4 U75B
-10 -8 18 0
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 16 0
1 U
3466 0 0
2
5.89983e-315 5.57017e-315
0
8 2-In OR~
219 1552 983 0 3 22
0 173 209 241
0
0 0 624 270
6 74LS32
-21 -24 21 -16
4 U75A
-10 -8 18 0
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 16 0
1 U
6910 0 0
2
5.89983e-315 5.5705e-315
0
8 2-In OR~
219 1324 981 0 3 22
0 178 214 246
0
0 0 624 270
6 74LS32
-21 -24 21 -16
4 U74D
-10 -8 18 0
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 15 0
1 U
8780 0 0
2
5.89983e-315 5.57082e-315
0
8 2-In OR~
219 1423 982 0 3 22
0 175 211 244
0
0 0 624 270
6 74LS32
-21 -24 21 -16
4 U74C
-10 -8 18 0
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 9 10 8 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 15 0
1 U
4905 0 0
2
5.89983e-315 5.57115e-315
0
8 2-In OR~
219 1390 982 0 3 22
0 176 212 243
0
0 0 624 270
6 74LS32
-21 -24 21 -16
4 U74B
-10 -8 18 0
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 15 0
1 U
3610 0 0
2
5.89983e-315 5.57147e-315
0
8 2-In OR~
219 1357 981 0 3 22
0 177 213 245
0
0 0 624 270
6 74LS32
-21 -24 21 -16
4 U74A
-10 -8 18 0
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 15 0
1 U
8414 0 0
2
5.89983e-315 5.57179e-315
0
8 2-In OR~
219 1514 588 0 3 22
0 182 218 250
0
0 0 624 270
6 74LS32
-21 -24 21 -16
4 U73D
-10 -8 18 0
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 14 0
1 U
5621 0 0
2
5.89983e-315 5.57212e-315
0
8 2-In OR~
219 1613 589 0 3 22
0 179 215 248
0
0 0 624 270
6 74LS32
-21 -24 21 -16
4 U73C
-10 -8 18 0
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 9 10 8 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 14 0
1 U
6801 0 0
2
5.89983e-315 5.57244e-315
0
8 2-In OR~
219 1580 589 0 3 22
0 180 216 247
0
0 0 624 270
6 74LS32
-21 -24 21 -16
4 U73B
-10 -8 18 0
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 14 0
1 U
8977 0 0
2
5.89983e-315 5.57276e-315
0
8 2-In OR~
219 1547 588 0 3 22
0 181 217 249
0
0 0 624 270
6 74LS32
-21 -24 21 -16
4 U73A
-10 -8 18 0
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 14 0
1 U
3646 0 0
2
5.89983e-315 5.57309e-315
0
8 2-In OR~
219 1315 589 0 3 22
0 186 222 254
0
0 0 624 270
6 74LS32
-21 -24 21 -16
4 U72D
-10 -8 18 0
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 13 0
1 U
7236 0 0
2
5.89983e-315 5.57341e-315
0
8 2-In OR~
219 1414 590 0 3 22
0 183 219 252
0
0 0 624 270
6 74LS32
-21 -24 21 -16
4 U72C
-10 -8 18 0
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 9 10 8 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 13 0
1 U
3586 0 0
2
5.89983e-315 5.57374e-315
0
8 2-In OR~
219 1381 590 0 3 22
0 184 220 251
0
0 0 624 270
6 74LS32
-21 -24 21 -16
4 U72B
-10 -8 18 0
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 13 0
1 U
4801 0 0
2
5.89983e-315 5.57406e-315
0
8 2-In OR~
219 1348 589 0 3 22
0 185 221 253
0
0 0 624 270
6 74LS32
-21 -24 21 -16
4 U72A
-10 -8 18 0
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 13 0
1 U
6689 0 0
2
5.89983e-315 5.57438e-315
0
8 2-In OR~
219 1541 186 0 3 22
0 189 225 52
0
0 0 624 270
6 74LS32
-21 -24 21 -16
4 U71D
-10 -8 18 0
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 12 0
1 U
7998 0 0
2
5.89983e-315 5.57471e-315
0
8 2-In OR~
219 1574 186 0 3 22
0 188 224 51
0
0 0 624 270
6 74LS32
-21 -24 21 -16
4 U71C
-10 -8 18 0
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 9 10 8 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 12 0
1 U
7254 0 0
2
5.89983e-315 5.57503e-315
0
8 2-In OR~
219 1607 186 0 3 22
0 187 223 50
0
0 0 624 270
6 74LS32
-21 -24 21 -16
4 U71B
-10 -8 18 0
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 12 0
1 U
6849 0 0
2
5.89983e-315 5.57535e-315
0
8 2-In OR~
219 1508 185 0 3 22
0 190 226 53
0
0 0 624 270
6 74LS32
-21 -24 21 -16
4 U71A
-10 -8 18 0
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 12 0
1 U
6684 0 0
2
5.89983e-315 5.57568e-315
0
8 2-In OR~
219 1311 182 0 3 22
0 194 230 57
0
0 0 624 270
6 74LS32
-21 -24 21 -16
4 U42D
-10 -8 18 0
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 11 0
1 U
3230 0 0
2
5.89983e-315 5.576e-315
0
8 2-In OR~
219 1410 184 0 3 22
0 191 227 54
0
0 0 624 270
6 74LS32
-21 -24 21 -16
4 U42C
-10 -8 18 0
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 9 10 8 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 11 0
1 U
5741 0 0
2
5.89983e-315 5.57633e-315
0
8 2-In OR~
219 1377 182 0 3 22
0 192 228 55
0
0 0 624 270
6 74LS32
-21 -24 21 -16
4 U42B
-10 -8 18 0
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 11 0
1 U
374 0 0
2
5.89983e-315 5.57665e-315
0
12 Quad D Flop~
47 2749 1430 0 9 19
0 255 256 257 258 262 261 260 259 162
0
0 0 4720 782
4 QDFF
-14 -44 14 -36
3 U67
-57 -4 -36 4
0
15 DVCC=16;DGND=8;
85 %D [%16bi %8bi %1i %2i %3i %4i %9i]
+ [%16bo %1o %2o %3o %4o %9o %5o %6o %7o %8o] %M
0
11 typeDigital
5 DIP16
19

0 1 2 3 4 5 6 7 8 9
1 2 3 4 5 6 7 8 9 0
65 0 0 0 1 0 0 0
1 U
5420 0 0
2
5.89983e-315 5.57697e-315
0
13 Quad 3-State~
48 2752 1484 0 9 19
0 262 261 260 259 190 189 188 187 7
0
0 0 4720 782
8 QUAD3STA
-28 -44 28 -36
3 U68
-60 -1 -39 7
0
15 DVCC=16;DGND=8;
85 %D [%16bi %8bi %1i %2i %3i %4i %9i]
+ [%16bo %1o %2o %3o %4o %9o %5o %6o %7o %8o] %M
0
12 type:digital
5 DIP16
19

0 1 2 3 4 5 6 7 8 9
1 2 3 4 5 6 7 8 9 0
65 0 0 0 1 0 0 0
1 U
8308 0 0
2
5.89983e-315 5.5773e-315
0
14 Logic Display~
6 2758 1360 0 1 2
10 258
0
0 0 53856 0
6 100MEG
3 -16 45 -8
3 L65
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
8158 0 0
2
5.89983e-315 5.57762e-315
0
14 Logic Display~
6 2725 1361 0 1 2
10 257
0
0 0 53856 0
6 100MEG
3 -16 45 -8
3 L66
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3979 0 0
2
5.89983e-315 5.57795e-315
0
14 Logic Display~
6 2694 1361 0 1 2
10 256
0
0 0 53856 0
6 100MEG
3 -16 45 -8
3 L67
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
9614 0 0
2
5.89983e-315 5.57827e-315
0
14 Logic Display~
6 2659 1361 0 1 2
10 255
0
0 0 53856 0
6 100MEG
3 -16 45 -8
3 L68
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
378 0 0
2
5.89983e-315 5.57859e-315
0
14 Logic Display~
6 2372 1369 0 1 2
10 263
0
0 0 53856 0
6 100MEG
3 -16 45 -8
3 L69
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
4325 0 0
2
5.89983e-315 5.57892e-315
0
14 Logic Display~
6 2407 1369 0 1 2
10 264
0
0 0 53856 0
6 100MEG
3 -16 45 -8
3 L70
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3282 0 0
2
5.89983e-315 5.57924e-315
0
14 Logic Display~
6 2438 1369 0 1 2
10 265
0
0 0 53856 0
6 100MEG
3 -16 45 -8
3 L71
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
5695 0 0
2
5.89983e-315 5.57956e-315
0
14 Logic Display~
6 2471 1368 0 1 2
10 266
0
0 0 53856 0
6 100MEG
3 -16 45 -8
3 L72
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3160 0 0
2
5.89983e-315 5.57989e-315
0
13 Quad 3-State~
48 2465 1492 0 9 19
0 270 269 268 267 194 193 192 191 7
0
0 0 4720 782
8 QUAD3STA
-28 -44 28 -36
3 U69
-60 -1 -39 7
0
15 DVCC=16;DGND=8;
85 %D [%16bi %8bi %1i %2i %3i %4i %9i]
+ [%16bo %1o %2o %3o %4o %9o %5o %6o %7o %8o] %M
0
12 type:digital
5 DIP16
19

0 1 2 3 4 5 6 7 8 9
1 2 3 4 5 6 7 8 9 0
65 0 0 0 1 0 0 0
1 U
5605 0 0
2
5.89983e-315 5.58021e-315
0
12 Quad D Flop~
47 2462 1438 0 9 19
0 263 264 265 266 270 269 268 267 162
0
0 0 4720 782
4 QDFF
-14 -44 14 -36
3 U70
-57 -4 -36 4
0
15 DVCC=16;DGND=8;
85 %D [%16bi %8bi %1i %2i %3i %4i %9i]
+ [%16bo %1o %2o %3o %4o %9o %5o %6o %7o %8o] %M
0
11 typeDigital
5 DIP16
19

0 1 2 3 4 5 6 7 8 9
1 2 3 4 5 6 7 8 9 0
65 0 0 0 1 0 0 0
1 U
8858 0 0
2
5.89983e-315 5.58054e-315
0
12 Quad D Flop~
47 2738 483 0 9 19
0 271 272 273 274 278 277 276 275 162
0
0 0 4720 782
4 QDFF
-14 -44 14 -36
3 U43
-57 -4 -36 4
0
15 DVCC=16;DGND=8;
85 %D [%16bi %8bi %1i %2i %3i %4i %9i]
+ [%16bo %1o %2o %3o %4o %9o %5o %6o %7o %8o] %M
0
11 typeDigital
5 DIP16
19

0 1 2 3 4 5 6 7 8 9
1 2 3 4 5 6 7 8 9 0
65 0 0 0 1 0 0 0
1 U
3697 0 0
2
5.89983e-315 5.58086e-315
0
13 Quad 3-State~
48 2741 537 0 9 19
0 278 277 276 275 218 217 216 215 8
0
0 0 4720 782
8 QUAD3STA
-28 -44 28 -36
3 U44
-60 -1 -39 7
0
15 DVCC=16;DGND=8;
85 %D [%16bi %8bi %1i %2i %3i %4i %9i]
+ [%16bo %1o %2o %3o %4o %9o %5o %6o %7o %8o] %M
0
12 type:digital
5 DIP16
19

0 1 2 3 4 5 6 7 8 9
1 2 3 4 5 6 7 8 9 0
65 0 0 0 1 0 0 0
1 U
4962 0 0
2
5.89983e-315 5.58118e-315
0
14 Logic Display~
6 2747 413 0 1 2
10 274
0
0 0 53856 0
6 100MEG
3 -16 45 -8
3 L17
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
6441 0 0
2
5.89983e-315 5.58151e-315
0
14 Logic Display~
6 2714 414 0 1 2
10 273
0
0 0 53856 0
6 100MEG
3 -16 45 -8
3 L18
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
4220 0 0
2
5.89983e-315 5.58183e-315
0
14 Logic Display~
6 2683 414 0 1 2
10 272
0
0 0 53856 0
6 100MEG
3 -16 45 -8
3 L19
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
9830 0 0
2
5.89983e-315 5.58215e-315
0
14 Logic Display~
6 2648 414 0 1 2
10 271
0
0 0 53856 0
6 100MEG
3 -16 45 -8
3 L20
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
7585 0 0
2
5.89983e-315 5.58248e-315
0
14 Logic Display~
6 2361 422 0 1 2
10 279
0
0 0 53856 0
6 100MEG
3 -16 45 -8
3 L21
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
5788 0 0
2
5.89983e-315 5.5828e-315
0
14 Logic Display~
6 2396 422 0 1 2
10 280
0
0 0 53856 0
6 100MEG
3 -16 45 -8
3 L22
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3262 0 0
2
5.89983e-315 5.58313e-315
0
14 Logic Display~
6 2427 422 0 1 2
10 281
0
0 0 53856 0
6 100MEG
3 -16 45 -8
3 L23
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
7575 0 0
2
5.89983e-315 5.58345e-315
0
14 Logic Display~
6 2460 421 0 1 2
10 282
0
0 0 53856 0
6 100MEG
3 -16 45 -8
3 L24
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
4232 0 0
2
5.89983e-315 5.58377e-315
0
13 Quad 3-State~
48 2454 545 0 9 19
0 286 285 284 283 222 221 220 219 8
0
0 0 4720 782
8 QUAD3STA
-28 -44 28 -36
3 U45
-60 -1 -39 7
0
15 DVCC=16;DGND=8;
85 %D [%16bi %8bi %1i %2i %3i %4i %9i]
+ [%16bo %1o %2o %3o %4o %9o %5o %6o %7o %8o] %M
0
12 type:digital
5 DIP16
19

0 1 2 3 4 5 6 7 8 9
1 2 3 4 5 6 7 8 9 0
65 0 0 0 1 0 0 0
1 U
8648 0 0
2
5.89983e-315 5.5841e-315
0
12 Quad D Flop~
47 2451 491 0 9 19
0 279 280 281 282 286 285 284 283 162
0
0 0 4720 782
4 QDFF
-14 -44 14 -36
3 U46
-57 -4 -36 4
0
15 DVCC=16;DGND=8;
85 %D [%16bi %8bi %1i %2i %3i %4i %9i]
+ [%16bo %1o %2o %3o %4o %9o %5o %6o %7o %8o] %M
0
11 typeDigital
5 DIP16
19

0 1 2 3 4 5 6 7 8 9
1 2 3 4 5 6 7 8 9 0
65 0 0 0 1 0 0 0
1 U
6524 0 0
2
5.89983e-315 5.58442e-315
0
7 Pulser~
4 2871 42 0 10 12
0 408 409 162 410 0 0 5 5 4
7
0
0 0 4656 0
0
3 V70
-10 -28 11 -20
0
0
0
0
0
4 SIP2
9

0 1 2 3 4 1 2 3 4 0
0 0 0 512 1 0 0 0
1 V
5265 0 0
2
5.89983e-315 5.58474e-315
0
12 Quad D Flop~
47 2753 1743 0 9 19
0 319 320 321 322 326 325 324 323 162
0
0 0 4720 782
4 QDFF
-14 -44 14 -36
3 U66
-57 -4 -36 4
0
15 DVCC=16;DGND=8;
85 %D [%16bi %8bi %1i %2i %3i %4i %9i]
+ [%16bo %1o %2o %3o %4o %9o %5o %6o %7o %8o] %M
0
11 typeDigital
5 DIP16
19

0 1 2 3 4 5 6 7 8 9
1 2 3 4 5 6 7 8 9 0
65 0 0 0 1 0 0 0
1 U
9322 0 0
2
5.89983e-315 5.58507e-315
0
13 Quad 3-State~
48 2756 1797 0 9 19
0 326 325 324 323 182 181 180 179 6
0
0 0 4720 782
8 QUAD3STA
-28 -44 28 -36
3 U65
-60 -1 -39 7
0
15 DVCC=16;DGND=8;
85 %D [%16bi %8bi %1i %2i %3i %4i %9i]
+ [%16bo %1o %2o %3o %4o %9o %5o %6o %7o %8o] %M
0
12 type:digital
5 DIP16
19

0 1 2 3 4 5 6 7 8 9
1 2 3 4 5 6 7 8 9 0
65 0 0 0 1 0 0 0
1 U
3103 0 0
2
5.89983e-315 5.58539e-315
0
14 Logic Display~
6 2762 1673 0 1 2
10 322
0
0 0 53856 0
6 100MEG
3 -16 45 -8
3 L64
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3156 0 0
2
5.89983e-315 5.58572e-315
0
14 Logic Display~
6 2729 1674 0 1 2
10 321
0
0 0 53856 0
6 100MEG
3 -16 45 -8
3 L63
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
7566 0 0
2
5.89983e-315 5.58604e-315
0
14 Logic Display~
6 2698 1674 0 1 2
10 320
0
0 0 53856 0
6 100MEG
3 -16 45 -8
3 L62
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3695 0 0
2
5.89983e-315 5.58636e-315
0
14 Logic Display~
6 2663 1674 0 1 2
10 319
0
0 0 53856 0
6 100MEG
3 -16 45 -8
3 L61
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
553 0 0
2
5.89983e-315 5.58669e-315
0
14 Logic Display~
6 2376 1682 0 1 2
10 327
0
0 0 53856 0
6 100MEG
3 -16 45 -8
3 L60
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
9168 0 0
2
5.89983e-315 5.58701e-315
0
14 Logic Display~
6 2411 1682 0 1 2
10 328
0
0 0 53856 0
6 100MEG
3 -16 45 -8
3 L59
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
869 0 0
2
5.89983e-315 5.58734e-315
0
14 Logic Display~
6 2442 1682 0 1 2
10 329
0
0 0 53856 0
6 100MEG
3 -16 45 -8
3 L58
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3125 0 0
2
5.89983e-315 5.58766e-315
0
14 Logic Display~
6 2475 1681 0 1 2
10 330
0
0 0 53856 0
6 100MEG
3 -16 45 -8
3 L57
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3845 0 0
2
5.89983e-315 5.58798e-315
0
13 Quad 3-State~
48 2469 1805 0 9 19
0 334 333 332 331 186 185 184 183 6
0
0 0 4720 782
8 QUAD3STA
-28 -44 28 -36
3 U64
-60 -1 -39 7
0
15 DVCC=16;DGND=8;
85 %D [%16bi %8bi %1i %2i %3i %4i %9i]
+ [%16bo %1o %2o %3o %4o %9o %5o %6o %7o %8o] %M
0
12 type:digital
5 DIP16
19

0 1 2 3 4 5 6 7 8 9
1 2 3 4 5 6 7 8 9 0
65 0 0 0 1 0 0 0
1 U
6597 0 0
2
5.89983e-315 5.58831e-315
0
12 Quad D Flop~
47 2466 1751 0 9 19
0 327 328 329 330 334 333 332 331 162
0
0 0 4720 782
4 QDFF
-14 -44 14 -36
3 U63
-57 -4 -36 4
0
15 DVCC=16;DGND=8;
85 %D [%16bi %8bi %1i %2i %3i %4i %9i]
+ [%16bo %1o %2o %3o %4o %9o %5o %6o %7o %8o] %M
0
11 typeDigital
5 DIP16
19

0 1 2 3 4 5 6 7 8 9
1 2 3 4 5 6 7 8 9 0
65 0 0 0 1 0 0 0
1 U
7163 0 0
2
5.89983e-315 5.58863e-315
0
12 Quad D Flop~
47 2750 2059 0 9 19
0 303 304 305 306 310 309 308 307 162
0
0 0 4720 782
4 QDFF
-14 -44 14 -36
3 U62
-57 -4 -36 4
0
15 DVCC=16;DGND=8;
85 %D [%16bi %8bi %1i %2i %3i %4i %9i]
+ [%16bo %1o %2o %3o %4o %9o %5o %6o %7o %8o] %M
0
11 typeDigital
5 DIP16
19

0 1 2 3 4 5 6 7 8 9
1 2 3 4 5 6 7 8 9 0
65 0 0 0 1 0 0 0
1 U
3127 0 0
2
5.89983e-315 5.58895e-315
0
13 Quad 3-State~
48 2753 2113 0 9 19
0 310 309 308 307 174 173 172 171 5
0
0 0 4720 782
8 QUAD3STA
-28 -44 28 -36
3 U61
-60 -1 -39 7
0
15 DVCC=16;DGND=8;
85 %D [%16bi %8bi %1i %2i %3i %4i %9i]
+ [%16bo %1o %2o %3o %4o %9o %5o %6o %7o %8o] %M
0
12 type:digital
5 DIP16
19

0 1 2 3 4 5 6 7 8 9
1 2 3 4 5 6 7 8 9 0
65 0 0 0 1 0 0 0
1 U
3815 0 0
2
5.89983e-315 5.58928e-315
0
14 Logic Display~
6 2759 1989 0 1 2
10 306
0
0 0 53856 0
6 100MEG
3 -16 45 -8
3 L56
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
9562 0 0
2
5.89983e-315 5.5896e-315
0
14 Logic Display~
6 2726 1990 0 1 2
10 305
0
0 0 53856 0
6 100MEG
3 -16 45 -8
3 L55
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
435 0 0
2
5.89983e-315 5.58993e-315
0
14 Logic Display~
6 2695 1990 0 1 2
10 304
0
0 0 53856 0
6 100MEG
3 -16 45 -8
3 L54
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
366 0 0
2
5.89983e-315 5.59025e-315
0
14 Logic Display~
6 2660 1990 0 1 2
10 303
0
0 0 53856 0
6 100MEG
3 -16 45 -8
3 L53
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
7315 0 0
2
5.89983e-315 5.59057e-315
0
14 Logic Display~
6 2373 1998 0 1 2
10 311
0
0 0 53856 0
6 100MEG
3 -16 45 -8
3 L52
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
328 0 0
2
5.89983e-315 5.5909e-315
0
14 Logic Display~
6 2408 1998 0 1 2
10 312
0
0 0 53856 0
6 100MEG
3 -16 45 -8
3 L51
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3936 0 0
2
5.89983e-315 5.59122e-315
0
14 Logic Display~
6 2439 1998 0 1 2
10 313
0
0 0 53856 0
6 100MEG
3 -16 45 -8
3 L50
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3965 0 0
2
5.89983e-315 5.59154e-315
0
14 Logic Display~
6 2472 1997 0 1 2
10 314
0
0 0 53856 0
6 100MEG
3 -16 45 -8
3 L49
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
4848 0 0
2
5.89983e-315 5.59187e-315
0
13 Quad 3-State~
48 2466 2121 0 9 19
0 318 317 316 315 178 177 176 175 5
0
0 0 4720 782
8 QUAD3STA
-28 -44 28 -36
3 U60
-60 -1 -39 7
0
15 DVCC=16;DGND=8;
85 %D [%16bi %8bi %1i %2i %3i %4i %9i]
+ [%16bo %1o %2o %3o %4o %9o %5o %6o %7o %8o] %M
0
12 type:digital
5 DIP16
19

0 1 2 3 4 5 6 7 8 9
1 2 3 4 5 6 7 8 9 0
65 0 0 0 1 0 0 0
1 U
859 0 0
2
5.89983e-315 5.59219e-315
0
12 Quad D Flop~
47 2463 2067 0 9 19
0 311 312 313 314 318 317 316 315 162
0
0 0 4720 782
4 QDFF
-14 -44 14 -36
3 U59
-57 -4 -36 4
0
15 DVCC=16;DGND=8;
85 %D [%16bi %8bi %1i %2i %3i %4i %9i]
+ [%16bo %1o %2o %3o %4o %9o %5o %6o %7o %8o] %M
0
11 typeDigital
5 DIP16
19

0 1 2 3 4 5 6 7 8 9
1 2 3 4 5 6 7 8 9 0
65 0 0 0 1 0 0 0
1 U
9385 0 0
2
5.89983e-315 5.59252e-315
0
12 Quad D Flop~
47 2751 2395 0 9 19
0 287 288 289 290 294 293 292 291 162
0
0 0 4720 782
4 QDFF
-14 -44 14 -36
3 U58
-57 -4 -36 4
0
15 DVCC=16;DGND=8;
85 %D [%16bi %8bi %1i %2i %3i %4i %9i]
+ [%16bo %1o %2o %3o %4o %9o %5o %6o %7o %8o] %M
0
11 typeDigital
5 DIP16
19

0 1 2 3 4 5 6 7 8 9
1 2 3 4 5 6 7 8 9 0
65 0 0 0 1 0 0 0
1 U
9823 0 0
2
5.89983e-315 5.59284e-315
0
13 Quad 3-State~
48 2754 2449 0 9 19
0 294 293 292 291 166 165 164 163 4
0
0 0 4720 782
8 QUAD3STA
-28 -44 28 -36
3 U57
-60 -1 -39 7
0
15 DVCC=16;DGND=8;
85 %D [%16bi %8bi %1i %2i %3i %4i %9i]
+ [%16bo %1o %2o %3o %4o %9o %5o %6o %7o %8o] %M
0
12 type:digital
5 DIP16
19

0 1 2 3 4 5 6 7 8 9
1 2 3 4 5 6 7 8 9 0
65 0 0 0 1 0 0 0
1 U
3509 0 0
2
5.89983e-315 5.59316e-315
0
14 Logic Display~
6 2760 2325 0 1 2
10 290
0
0 0 53856 0
6 100MEG
3 -16 45 -8
3 L48
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
7783 0 0
2
5.89983e-315 5.59349e-315
0
14 Logic Display~
6 2727 2326 0 1 2
10 289
0
0 0 53856 0
6 100MEG
3 -16 45 -8
3 L47
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
9834 0 0
2
5.89983e-315 5.59381e-315
0
14 Logic Display~
6 2696 2326 0 1 2
10 288
0
0 0 53856 0
6 100MEG
3 -16 45 -8
3 L46
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
4814 0 0
2
5.89983e-315 5.59413e-315
0
14 Logic Display~
6 2661 2326 0 1 2
10 287
0
0 0 53856 0
6 100MEG
3 -16 45 -8
3 L45
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3513 0 0
2
5.89983e-315 5.59446e-315
0
14 Logic Display~
6 2374 2334 0 1 2
10 295
0
0 0 53856 0
6 100MEG
3 -16 45 -8
3 L44
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
7249 0 0
2
5.89983e-315 5.59478e-315
0
14 Logic Display~
6 2409 2334 0 1 2
10 296
0
0 0 53856 0
6 100MEG
3 -16 45 -8
3 L43
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
8268 0 0
2
5.89983e-315 5.59511e-315
0
14 Logic Display~
6 2440 2334 0 1 2
10 297
0
0 0 53856 0
6 100MEG
3 -16 45 -8
3 L42
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
8799 0 0
2
5.89983e-315 5.59527e-315
0
14 Logic Display~
6 2473 2333 0 1 2
10 298
0
0 0 53856 0
6 100MEG
3 -16 45 -8
3 L41
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3830 0 0
2
5.89983e-315 5.59543e-315
0
13 Quad 3-State~
48 2467 2457 0 9 19
0 302 301 300 299 170 169 168 167 4
0
0 0 4720 782
8 QUAD3STA
-28 -44 28 -36
3 U56
-60 -1 -39 7
0
15 DVCC=16;DGND=8;
85 %D [%16bi %8bi %1i %2i %3i %4i %9i]
+ [%16bo %1o %2o %3o %4o %9o %5o %6o %7o %8o] %M
0
12 type:digital
5 DIP16
19

0 1 2 3 4 5 6 7 8 9
1 2 3 4 5 6 7 8 9 0
65 0 0 0 1 0 0 0
1 U
8985 0 0
2
5.89983e-315 5.59559e-315
0
12 Quad D Flop~
47 2464 2403 0 9 19
0 295 296 297 298 302 301 300 299 162
0
0 0 4720 782
4 QDFF
-14 -44 14 -36
3 U55
-57 -4 -36 4
0
15 DVCC=16;DGND=8;
85 %D [%16bi %8bi %1i %2i %3i %4i %9i]
+ [%16bo %1o %2o %3o %4o %9o %5o %6o %7o %8o] %M
0
11 typeDigital
5 DIP16
19

0 1 2 3 4 5 6 7 8 9
1 2 3 4 5 6 7 8 9 0
65 0 0 0 1 0 0 0
1 U
3678 0 0
2
5.89983e-315 5.59575e-315
0
12 Quad D Flop~
47 2456 1129 0 9 19
0 343 344 345 346 206 205 204 203 162
0
0 0 4720 782
4 QDFF
-14 -44 14 -36
3 U54
-57 -4 -36 4
0
15 DVCC=16;DGND=8;
85 %D [%16bi %8bi %1i %2i %3i %4i %9i]
+ [%16bo %1o %2o %3o %4o %9o %5o %6o %7o %8o] %M
0
11 typeDigital
5 DIP16
19

0 1 2 3 4 5 6 7 8 9
1 2 3 4 5 6 7 8 9 0
65 0 0 0 1 0 0 0
1 U
3939 0 0
2
5.89983e-315 5.59592e-315
0
13 Quad 3-State~
48 2459 1183 0 9 19
0 206 205 204 203 202 201 200 199 105
0
0 0 4720 782
8 QUAD3STA
-28 -44 28 -36
3 U53
-64 -1 -43 7
0
15 DVCC=16;DGND=8;
85 %D [%16bi %8bi %1i %2i %3i %4i %9i]
+ [%16bo %1o %2o %3o %4o %9o %5o %6o %7o %8o] %M
0
12 type:digital
5 DIP16
19

0 1 2 3 4 5 6 7 8 9
1 2 3 4 5 6 7 8 9 0
65 0 0 0 1 0 0 0
1 U
8325 0 0
2
5.89983e-315 5.59608e-315
0
14 Logic Display~
6 2465 1059 0 1 2
10 346
0
0 0 53856 0
6 100MEG
3 -16 45 -8
3 L40
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
7461 0 0
2
5.89983e-315 5.59624e-315
0
14 Logic Display~
6 2432 1060 0 1 2
10 345
0
0 0 53856 0
6 100MEG
3 -16 45 -8
3 L39
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
7656 0 0
2
5.89983e-315 5.5964e-315
0
14 Logic Display~
6 2401 1060 0 1 2
10 344
0
0 0 53856 0
6 100MEG
3 -16 45 -8
3 L38
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3602 0 0
2
5.89983e-315 5.59656e-315
0
14 Logic Display~
6 2366 1060 0 1 2
10 343
0
0 0 53856 0
6 100MEG
3 -16 45 -8
3 L37
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3383 0 0
2
5.89983e-315 5.59673e-315
0
14 Logic Display~
6 2653 1052 0 1 2
10 335
0
0 0 53856 0
6 100MEG
3 -16 45 -8
3 L36
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3845 0 0
2
5.89983e-315 5.59689e-315
0
14 Logic Display~
6 2688 1052 0 1 2
10 336
0
0 0 53856 0
6 100MEG
3 -16 45 -8
3 L35
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
571 0 0
2
5.89983e-315 5.59705e-315
0
14 Logic Display~
6 2719 1052 0 1 2
10 337
0
0 0 53856 0
6 100MEG
3 -16 45 -8
3 L34
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3172 0 0
2
5.89983e-315 5.59721e-315
0
14 Logic Display~
6 2752 1051 0 1 2
10 338
0
0 0 53856 0
6 100MEG
3 -16 45 -8
3 L33
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3250 0 0
2
5.89983e-315 5.59737e-315
0
13 Quad 3-State~
48 2746 1175 0 9 19
0 342 341 340 339 198 197 196 195 105
0
0 0 4720 782
8 QUAD3STA
-28 -44 28 -36
3 U52
-60 -1 -39 7
0
15 DVCC=16;DGND=8;
85 %D [%16bi %8bi %1i %2i %3i %4i %9i]
+ [%16bo %1o %2o %3o %4o %9o %5o %6o %7o %8o] %M
0
12 type:digital
5 DIP16
19

0 1 2 3 4 5 6 7 8 9
1 2 3 4 5 6 7 8 9 0
65 0 0 0 1 0 0 0
1 U
3865 0 0
2
5.89983e-315 5.59753e-315
0
12 Quad D Flop~
47 2743 1121 0 9 19
0 335 336 337 338 342 341 340 339 162
0
0 0 4720 782
4 QDFF
-14 -44 14 -36
3 U51
-57 -4 -36 4
0
15 DVCC=16;DGND=8;
85 %D [%16bi %8bi %1i %2i %3i %4i %9i]
+ [%16bo %1o %2o %3o %4o %9o %5o %6o %7o %8o] %M
0
11 typeDigital
5 DIP16
19

0 1 2 3 4 5 6 7 8 9
1 2 3 4 5 6 7 8 9 0
65 0 0 0 1 0 0 0
1 U
3253 0 0
2
5.89983e-315 5.5977e-315
0
12 Quad D Flop~
47 2455 793 0 9 19
0 355 356 357 358 362 361 360 359 162
0
0 0 4720 782
4 QDFF
-14 -44 14 -36
3 U50
-57 -4 -36 4
0
15 DVCC=16;DGND=8;
85 %D [%16bi %8bi %1i %2i %3i %4i %9i]
+ [%16bo %1o %2o %3o %4o %9o %5o %6o %7o %8o] %M
0
11 typeDigital
5 DIP16
19

0 1 2 3 4 5 6 7 8 9
1 2 3 4 5 6 7 8 9 0
65 0 0 0 1 0 0 0
1 U
6957 0 0
2
5.89983e-315 5.59786e-315
0
13 Quad 3-State~
48 2458 847 0 9 19
0 362 361 360 359 214 213 212 211 108
0
0 0 4720 782
8 QUAD3STA
-28 -44 28 -36
3 U49
-60 -1 -39 7
0
15 DVCC=16;DGND=8;
85 %D [%16bi %8bi %1i %2i %3i %4i %9i]
+ [%16bo %1o %2o %3o %4o %9o %5o %6o %7o %8o] %M
0
12 type:digital
5 DIP16
19

0 1 2 3 4 5 6 7 8 9
1 2 3 4 5 6 7 8 9 0
65 0 0 0 1 0 0 0
1 U
9668 0 0
2
5.89983e-315 5.59802e-315
0
14 Logic Display~
6 2464 723 0 1 2
10 358
0
0 0 53856 0
6 100MEG
3 -16 45 -8
3 L32
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3765 0 0
2
5.89983e-315 5.59818e-315
0
14 Logic Display~
6 2431 724 0 1 2
10 357
0
0 0 53856 0
6 100MEG
3 -16 45 -8
3 L31
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
4286 0 0
2
5.89983e-315 5.59834e-315
0
14 Logic Display~
6 2400 724 0 1 2
10 356
0
0 0 53856 0
6 100MEG
3 -16 45 -8
3 L30
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
76 0 0
2
5.89983e-315 5.59851e-315
0
14 Logic Display~
6 2365 724 0 1 2
10 355
0
0 0 53856 0
6 100MEG
3 -16 45 -8
3 L29
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
9206 0 0
2
5.89983e-315 5.59867e-315
0
14 Logic Display~
6 2652 716 0 1 2
10 347
0
0 0 53856 0
6 100MEG
3 -16 45 -8
3 L28
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
9169 0 0
2
5.89983e-315 5.59883e-315
0
14 Logic Display~
6 2687 716 0 1 2
10 348
0
0 0 53856 0
6 100MEG
3 -16 45 -8
3 L27
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
9384 0 0
2
5.89983e-315 5.59899e-315
0
14 Logic Display~
6 2718 716 0 1 2
10 349
0
0 0 53856 0
6 100MEG
3 -16 45 -8
3 L26
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
6605 0 0
2
5.89983e-315 5.59915e-315
0
14 Logic Display~
6 2751 715 0 1 2
10 350
0
0 0 53856 0
6 100MEG
3 -16 45 -8
3 L25
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3294 0 0
2
5.89983e-315 5.59932e-315
0
13 Quad 3-State~
48 2745 839 0 9 19
0 354 353 352 351 210 209 208 207 108
0
0 0 4720 782
8 QUAD3STA
-28 -44 28 -36
3 U48
-60 -1 -39 7
0
15 DVCC=16;DGND=8;
85 %D [%16bi %8bi %1i %2i %3i %4i %9i]
+ [%16bo %1o %2o %3o %4o %9o %5o %6o %7o %8o] %M
0
12 type:digital
5 DIP16
19

0 1 2 3 4 5 6 7 8 9
1 2 3 4 5 6 7 8 9 0
65 0 0 0 1 0 0 0
1 U
633 0 0
2
5.89983e-315 5.59948e-315
0
12 Quad D Flop~
47 2742 785 0 9 19
0 347 348 349 350 354 353 352 351 162
0
0 0 4720 782
4 QDFF
-14 -44 14 -36
3 U47
-57 -4 -36 4
0
15 DVCC=16;DGND=8;
85 %D [%16bi %8bi %1i %2i %3i %4i %9i]
+ [%16bo %1o %2o %3o %4o %9o %5o %6o %7o %8o] %M
0
11 typeDigital
5 DIP16
19

0 1 2 3 4 5 6 7 8 9
1 2 3 4 5 6 7 8 9 0
65 0 0 0 1 0 0 0
1 U
3179 0 0
2
5.89983e-315 5.59964e-315
0
12 Quad D Flop~
47 2735 202 0 9 19
0 363 364 365 366 370 369 368 367 162
0
0 0 4720 782
4 QDFF
-14 -44 14 -36
3 U37
-57 -4 -36 4
0
15 DVCC=16;DGND=8;
85 %D [%16bi %8bi %1i %2i %3i %4i %9i]
+ [%16bo %1o %2o %3o %4o %9o %5o %6o %7o %8o] %M
0
11 typeDigital
5 DIP16
19

0 1 2 3 4 5 6 7 8 9
1 2 3 4 5 6 7 8 9 0
65 0 0 0 1 0 0 0
1 U
3900 0 0
2
5.89983e-315 5.5998e-315
0
13 Quad 3-State~
48 2738 256 0 9 19
0 370 369 368 367 226 225 224 223 60
0
0 0 4720 782
8 QUAD3STA
-28 -44 28 -36
3 U36
-60 -1 -39 7
0
15 DVCC=16;DGND=8;
85 %D [%16bi %8bi %1i %2i %3i %4i %9i]
+ [%16bo %1o %2o %3o %4o %9o %5o %6o %7o %8o] %M
0
12 type:digital
5 DIP16
19

0 1 2 3 4 5 6 7 8 9
1 2 3 4 5 6 7 8 9 0
65 0 0 0 1 0 0 0
1 U
8562 0 0
2
5.89983e-315 5.59996e-315
0
14 Logic Display~
6 2744 132 0 1 2
10 366
0
0 0 53856 0
6 100MEG
3 -16 45 -8
3 L16
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3117 0 0
2
5.89983e-315 5.60012e-315
0
14 Logic Display~
6 2711 133 0 1 2
10 365
0
0 0 53856 0
6 100MEG
3 -16 45 -8
3 L15
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3703 0 0
2
5.89983e-315 5.60029e-315
0
14 Logic Display~
6 2680 133 0 1 2
10 364
0
0 0 53856 0
6 100MEG
3 -16 45 -8
3 L14
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
9799 0 0
2
5.89983e-315 5.60045e-315
0
14 Logic Display~
6 2645 133 0 1 2
10 363
0
0 0 53856 0
6 100MEG
3 -16 45 -8
3 L13
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
668 0 0
2
5.89983e-315 5.60061e-315
0
14 Logic Display~
6 2358 141 0 1 2
10 371
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L9
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3928 0 0
2
5.89983e-315 5.60077e-315
0
14 Logic Display~
6 2393 141 0 1 2
10 372
0
0 0 53856 0
6 100MEG
3 -16 45 -8
3 L10
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
378 0 0
2
5.89983e-315 5.60093e-315
0
14 Logic Display~
6 2424 141 0 1 2
10 373
0
0 0 53856 0
6 100MEG
3 -16 45 -8
3 L11
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3579 0 0
2
5.89983e-315 5.6011e-315
0
14 Logic Display~
6 2457 140 0 1 2
10 374
0
0 0 53856 0
6 100MEG
3 -16 45 -8
3 L12
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
9637 0 0
2
5.89983e-315 5.60126e-315
0
8 2-In OR~
219 1344 182 0 3 22
0 193 229 56
0
0 0 624 270
6 74LS32
-21 -24 21 -16
4 U42A
-10 -8 18 0
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 11 0
1 U
6196 0 0
2
5.89983e-315 5.60142e-315
0
13 Quad 3-State~
48 2451 264 0 9 19
0 379 378 377 376 230 229 228 227 60
0
0 0 4720 782
8 QUAD3STA
-28 -44 28 -36
3 U41
-60 -1 -39 7
0
15 DVCC=16;DGND=8;
85 %D [%16bi %8bi %1i %2i %3i %4i %9i]
+ [%16bo %1o %2o %3o %4o %9o %5o %6o %7o %8o] %M
0
12 type:digital
5 DIP16
19

0 1 2 3 4 5 6 7 8 9
1 2 3 4 5 6 7 8 9 0
65 0 0 0 1 0 0 0
1 U
6292 0 0
2
5.89983e-315 5.60158e-315
0
12 Quad D Flop~
47 2448 210 0 9 19
0 371 372 373 374 379 378 377 376 162
0
0 0 4720 782
4 QDFF
-14 -44 14 -36
3 U40
-57 -4 -36 4
0
15 DVCC=16;DGND=8;
85 %D [%16bi %8bi %1i %2i %3i %4i %9i]
+ [%16bo %1o %2o %3o %4o %9o %5o %6o %7o %8o] %M
0
11 typeDigital
5 DIP16
19

0 1 2 3 4 5 6 7 8 9
1 2 3 4 5 6 7 8 9 0
65 0 0 0 1 0 0 0
1 U
3605 0 0
2
5.89983e-315 5.60174e-315
0
14 Logic Display~
6 486 595 0 1 2
10 380
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L8
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3697 0 0
2
44331.3 33
0
14 Logic Display~
6 487 538 0 1 2
10 3
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L7
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3620 0 0
2
44331.3 34
0
9 Inverter~
13 193 369 0 2 22
0 384 383
0
0 0 624 0
6 74LS04
-21 -19 21 -11
3 U3D
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 9 8 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 4 1 0
1 U
8890 0 0
2
44331.3 35
0
14 Logic Display~
6 163 350 0 1 2
10 384
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L6
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
8729 0 0
2
44331.3 36
0
13 Quad 3-State~
48 247 486 0 9 19
0 388 389 390 391 381 380 3 382 383
0
0 0 4720 692
8 QUAD3STA
-28 -44 28 -36
3 U38
-11 46 10 54
0
15 DVCC=16;DGND=8;
85 %D [%16bi %8bi %1i %2i %3i %4i %9i]
+ [%16bo %1o %2o %3o %4o %9o %5o %6o %7o %8o] %M
0
12 type:digital
5 DIP16
19

0 1 2 3 4 5 6 7 8 9
1 2 3 4 5 6 7 8 9 0
65 0 0 0 1 0 0 0
1 U
47 0 0
2
44331.3 37
0
8 4-In OR~
219 1480 2016 0 5 22
0 385 386 387 375 41
0
0 0 624 0
4 4072
-14 -24 14 -16
4 U39A
-6 -25 22 -17
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
12 type:digital
5 DIP14
22

0 2 3 4 5 1 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 0 2 1 10 0
1 U
4533 0 0
2
44331.3 38
0
14 Logic Display~
6 181 453 0 1 2
10 390
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L3
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
9356 0 0
2
44331.3 39
0
14 Logic Display~
6 196 453 0 1 2
10 389
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L4
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3206 0 0
2
44331.3 40
0
14 Logic Display~
6 211 453 0 1 2
10 388
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L5
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
9695 0 0
2
44331.3 41
0
14 Logic Display~
6 165 453 0 1 2
10 391
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L2
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
5663 0 0
2
44331.3 42
0
4 4514
219 1621 2039 0 30 45
0 382 3 380 381 41 411 155 154 153
152 151 150 147 146 145 144 143 142 141
140 139 138 0 0 0 0 0 0 0
5
0
0 0 4848 692
4 4514
-14 -87 14 -79
2 U6
-7 -88 7 -80
0
16 DVDD=24;DGND=12;
155 %D [%24bi %12bi %1i %2i %3i %4i %5i %6i]
+ [%24bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o %15o %16o %17o %18o %19o %20o %21o %22o] %M
0
12 type:digital
5 DIP24
45

0 22 21 3 2 1 23 11 9 10
8 7 6 5 4 18 17 20 19 14
13 16 15 22 21 3 2 1 23 11
9 10 8 7 6 5 4 18 17 20
19 14 13 16 15 0
65 0 0 512 1 0 0 0
1 U
3199 0 0
2
44331.3 43
0
12 D Flip-Flop~
219 1108 1639 0 4 9
0 119 118 412 96
0
0 0 4720 0
3 DFF
-10 -53 11 -45
3 U34
-11 -55 10 -47
0
14 DVCC=6;DGND=5;
47 %D [%6bi %5bi %1i %2i][%6bo %1o %2o %3o %4o] %M
0
11 typeDigital
4 DIP6
9

0 1 2 3 4 1 2 3 4 0
65 0 0 512 1 0 0 0
1 U
7900 0 0
2
44331.3 44
0
12 D Flip-Flop~
219 949 1642 0 4 9
0 128 127 413 97
0
0 0 4720 0
3 DFF
-10 -53 11 -45
3 U35
-11 -55 10 -47
0
14 DVCC=6;DGND=5;
47 %D [%6bi %5bi %1i %2i][%6bo %1o %2o %3o %4o] %M
0
11 typeDigital
4 DIP6
9

0 1 2 3 4 1 2 3 4 0
65 0 0 512 1 0 0 0
1 U
7793 0 0
2
44331.3 45
0
9 2-In AND~
219 1250 1695 0 3 22
0 97 375 95
0
0 0 624 0
6 74LS08
-21 -24 21 -16
4 U20C
-13 -9 15 -1
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 8 0
1 U
3190 0 0
2
44331.3 46
0
6 74266~
219 1166 1738 0 3 22
0 96 382 375
0
0 0 624 0
7 74LS266
-24 -24 25 -16
4 U11D
-3 -12 25 -4
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 6 0
1 U
8930 0 0
2
44331.3 47
0
13 Quad 3-State~
48 1397 1686 0 9 19
0 28 27 26 25 70 69 68 67 394
0
0 0 4720 782
8 QUAD3STA
-28 -44 28 -36
3 U32
-60 -1 -39 7
0
15 DVCC=16;DGND=8;
85 %D [%16bi %8bi %1i %2i %3i %4i %9i]
+ [%16bo %1o %2o %3o %4o %9o %5o %6o %7o %8o] %M
0
12 type:digital
5 DIP16
19

0 1 2 3 4 5 6 7 8 9
1 2 3 4 5 6 7 8 9 0
65 0 0 0 1 0 0 0
1 U
9797 0 0
2
44331.3 48
0
12 Quad D Flop~
47 1394 1570 0 9 19
0 238 237 235 236 28 27 26 25 149
0
0 0 4720 782
4 QDFF
-14 -44 14 -36
3 U33
-57 -4 -36 4
0
15 DVCC=16;DGND=8;
85 %D [%16bi %8bi %1i %2i %3i %4i %9i]
+ [%16bo %1o %2o %3o %4o %9o %5o %6o %7o %8o] %M
0
11 typeDigital
5 DIP16
19

0 1 2 3 4 5 6 7 8 9
1 2 3 4 5 6 7 8 9 0
65 0 0 0 1 0 0 0
1 U
3472 0 0
2
44331.3 49
0
5 7412~
219 1318 1780 0 4 22
0 95 393 392 394
0
0 0 624 0
4 7412
-7 -24 21 -16
4 U29B
-14 -9 14 -1
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 1 2 8 9 3 4 5 6 1
2 8 9 11 12 13 10 0 0 0
0 6 0
65 0 0 0 3 2 9 0
1 U
4304 0 0
2
44331.3 50
0
5 7412~
219 1398 1829 0 4 22
0 95 393 381 395
0
0 0 624 0
4 7412
-7 -24 21 -16
4 U29A
-13 -13 15 -5
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 3 4 5 6 3 4 5 6 1
2 8 9 11 12 13 10 0 0 0
0 6 0
65 0 0 0 3 1 9 0
1 U
9362 0 0
2
44331.3 51
0
12 Quad D Flop~
47 1584 1573 0 9 19
0 234 233 231 232 12 11 10 9 148
0
0 0 4720 782
4 QDFF
-14 -44 14 -36
3 U30
-57 -4 -36 4
0
15 DVCC=16;DGND=8;
85 %D [%16bi %8bi %1i %2i %3i %4i %9i]
+ [%16bo %1o %2o %3o %4o %9o %5o %6o %7o %8o] %M
0
11 typeDigital
5 DIP16
19

0 1 2 3 4 5 6 7 8 9
1 2 3 4 5 6 7 8 9 0
65 0 0 0 1 0 0 0
1 U
8808 0 0
2
44331.3 52
0
13 Quad 3-State~
48 1587 1686 0 9 19
0 12 11 10 9 66 65 64 63 395
0
0 0 4720 782
8 QUAD3STA
-28 -44 28 -36
3 U31
-60 -1 -39 7
0
15 DVCC=16;DGND=8;
85 %D [%16bi %8bi %1i %2i %3i %4i %9i]
+ [%16bo %1o %2o %3o %4o %9o %5o %6o %7o %8o] %M
0
12 type:digital
5 DIP16
19

0 1 2 3 4 5 6 7 8 9
1 2 3 4 5 6 7 8 9 0
65 0 0 0 1 0 0 0
1 U
3972 0 0
2
44331.3 53
0
12 D Flip-Flop~
219 1108 1109 0 4 9
0 121 120 414 100
0
0 0 4720 0
3 DFF
-10 -53 11 -45
3 U28
-11 -55 10 -47
0
14 DVCC=6;DGND=5;
47 %D [%6bi %5bi %1i %2i][%6bo %1o %2o %3o %4o] %M
0
11 typeDigital
4 DIP6
9

0 1 2 3 4 1 2 3 4 0
65 0 0 512 1 0 0 0
1 U
3869 0 0
2
44331.3 54
0
12 D Flip-Flop~
219 937 1106 0 4 9
0 131 130 415 99
0
0 0 4720 0
3 DFF
-10 -53 11 -45
3 U27
-11 -55 10 -47
0
14 DVCC=6;DGND=5;
47 %D [%6bi %5bi %1i %2i][%6bo %1o %2o %3o %4o] %M
0
11 typeDigital
4 DIP6
9

0 1 2 3 4 1 2 3 4 0
65 0 0 512 1 0 0 0
1 U
9376 0 0
2
44331.3 55
0
9 2-In AND~
219 1238 1140 0 3 22
0 99 387 98
0
0 0 624 0
6 74LS08
-21 -24 21 -16
4 U20B
-12 -9 16 -1
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 8 0
1 U
8287 0 0
2
44331.3 56
0
6 74266~
219 1163 1183 0 3 22
0 100 382 387
0
0 0 624 0
7 74LS266
-24 -24 25 -16
4 U11C
-3 -12 25 -4
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 8 9 10 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 6 0
1 U
342 0 0
2
44331.3 57
0
13 Quad 3-State~
48 1390 1154 0 9 19
0 32 31 30 29 78 77 76 75 397
0
0 0 4720 782
8 QUAD3STA
-28 -44 28 -36
3 U26
-60 -1 -39 7
0
15 DVCC=16;DGND=8;
85 %D [%16bi %8bi %1i %2i %3i %4i %9i]
+ [%16bo %1o %2o %3o %4o %9o %5o %6o %7o %8o] %M
0
12 type:digital
5 DIP16
19

0 1 2 3 4 5 6 7 8 9
1 2 3 4 5 6 7 8 9 0
65 0 0 0 1 0 0 0
1 U
4378 0 0
2
44331.3 58
0
12 Quad D Flop~
47 1387 1050 0 9 19
0 246 245 243 244 32 31 30 29 157
0
0 0 4720 782
4 QDFF
-14 -44 14 -36
3 U24
-57 -4 -36 4
0
15 DVCC=16;DGND=8;
85 %D [%16bi %8bi %1i %2i %3i %4i %9i]
+ [%16bo %1o %2o %3o %4o %9o %5o %6o %7o %8o] %M
0
11 typeDigital
5 DIP16
19

0 1 2 3 4 5 6 7 8 9
1 2 3 4 5 6 7 8 9 0
65 0 0 0 1 0 0 0
1 U
6617 0 0
2
44331.3 59
0
5 7412~
219 1304 1227 0 4 22
0 98 396 392 397
0
0 0 624 0
4 7412
-7 -24 21 -16
4 U15C
-14 -9 14 -1
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 11 12 13 10 3 4 5 6 1
2 8 9 11 12 13 10 0 0 0
0 6 0
65 0 0 0 3 3 7 0
1 U
6432 0 0
2
44331.3 60
0
5 7412~
219 1393 1287 0 4 22
0 98 396 381 398
0
0 0 624 0
4 7412
-7 -24 21 -16
4 U15B
-13 -13 15 -5
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 1 2 8 9 3 4 5 6 1
2 8 9 11 12 13 10 0 0 0
0 6 0
65 0 0 0 3 2 7 0
1 U
6470 0 0
2
44331.3 61
0
12 Quad D Flop~
47 1582 1056 0 9 19
0 242 241 239 240 16 15 14 13 156
0
0 0 4720 782
4 QDFF
-14 -44 14 -36
3 U23
-57 -4 -36 4
0
15 DVCC=16;DGND=8;
85 %D [%16bi %8bi %1i %2i %3i %4i %9i]
+ [%16bo %1o %2o %3o %4o %9o %5o %6o %7o %8o] %M
0
11 typeDigital
5 DIP16
19

0 1 2 3 4 5 6 7 8 9
1 2 3 4 5 6 7 8 9 0
65 0 0 0 1 0 0 0
1 U
3215 0 0
2
44331.3 62
0
13 Quad 3-State~
48 1585 1156 0 9 19
0 16 15 14 13 74 73 72 71 398
0
0 0 4720 782
8 QUAD3STA
-28 -44 28 -36
3 U22
-60 -1 -39 7
0
15 DVCC=16;DGND=8;
85 %D [%16bi %8bi %1i %2i %3i %4i %9i]
+ [%16bo %1o %2o %3o %4o %9o %5o %6o %7o %8o] %M
0
12 type:digital
5 DIP16
19

0 1 2 3 4 5 6 7 8 9
1 2 3 4 5 6 7 8 9 0
65 0 0 0 1 0 0 0
1 U
8677 0 0
2
44331.3 63
0
6 74266~
219 1141 790 0 3 22
0 102 382 386
0
0 0 624 0
7 74LS266
-24 -24 25 -16
4 U11B
-3 -12 25 -4
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 5 6 4 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 6 0
1 U
8201 0 0
2
44331.3 64
0
9 2-In AND~
219 1216 758 0 3 22
0 61 386 101
0
0 0 624 0
6 74LS08
-21 -24 21 -16
4 U20A
-12 -12 16 -4
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 8 0
1 U
4920 0 0
2
44331.3 65
0
12 D Flip-Flop~
219 915 729 0 4 9
0 134 133 416 61
0
0 0 4720 0
3 DFF
-10 -53 11 -45
3 U19
-11 -55 10 -47
0
14 DVCC=6;DGND=5;
47 %D [%6bi %5bi %1i %2i][%6bo %1o %2o %3o %4o] %M
0
11 typeDigital
4 DIP6
9

0 1 2 3 4 1 2 3 4 0
65 0 0 512 1 0 0 0
1 U
911 0 0
2
44331.3 66
0
12 D Flip-Flop~
219 1084 732 0 4 9
0 123 122 417 102
0
0 0 4720 0
3 DFF
-10 -53 11 -45
3 U18
-11 -55 10 -47
0
14 DVCC=6;DGND=5;
47 %D [%6bi %5bi %1i %2i][%6bo %1o %2o %3o %4o] %M
0
11 typeDigital
4 DIP6
9

0 1 2 3 4 1 2 3 4 0
65 0 0 512 1 0 0 0
1 U
4377 0 0
2
44331.3 67
0
5 7412~
219 1293 838 0 4 22
0 101 399 392 401
0
0 0 624 0
4 7412
-7 -24 21 -16
3 U9C
-11 -12 10 -4
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 11 12 13 10 3 4 5 6 1
2 8 9 11 12 13 10 0 0 0
0 6 0
65 0 0 0 3 3 4 0
1 U
3916 0 0
2
44331.3 68
0
12 Quad D Flop~
47 1378 662 0 9 19
0 254 253 251 252 36 35 34 33 159
0
0 0 4720 782
4 QDFF
-14 -44 14 -36
3 U13
-57 -4 -36 4
0
15 DVCC=16;DGND=8;
85 %D [%16bi %8bi %1i %2i %3i %4i %9i]
+ [%16bo %1o %2o %3o %4o %9o %5o %6o %7o %8o] %M
0
11 typeDigital
5 DIP16
19

0 1 2 3 4 5 6 7 8 9
1 2 3 4 5 6 7 8 9 0
65 0 0 0 1 0 0 0
1 U
4666 0 0
2
44331.3 69
0
13 Quad 3-State~
48 1381 747 0 9 19
0 36 35 34 33 94 93 92 91 401
0
0 0 4720 782
8 QUAD3STA
-28 -44 28 -36
3 U14
-60 -1 -39 7
0
15 DVCC=16;DGND=8;
85 %D [%16bi %8bi %1i %2i %3i %4i %9i]
+ [%16bo %1o %2o %3o %4o %9o %5o %6o %7o %8o] %M
0
12 type:digital
5 DIP16
19

0 1 2 3 4 5 6 7 8 9
1 2 3 4 5 6 7 8 9 0
65 0 0 0 1 0 0 0
1 U
7507 0 0
2
44331.3 70
0
13 Quad 3-State~
48 1580 748 0 9 19
0 20 19 18 17 82 81 80 79 402
0
0 0 4720 782
8 QUAD3STA
-28 -44 28 -36
3 U17
-60 -1 -39 7
0
15 DVCC=16;DGND=8;
85 %D [%16bi %8bi %1i %2i %3i %4i %9i]
+ [%16bo %1o %2o %3o %4o %9o %5o %6o %7o %8o] %M
0
12 type:digital
5 DIP16
19

0 1 2 3 4 5 6 7 8 9
1 2 3 4 5 6 7 8 9 0
65 0 0 0 1 0 0 0
1 U
4350 0 0
2
44331.3 71
0
12 Quad D Flop~
47 1577 661 0 9 19
0 250 249 247 248 20 19 18 17 158
0
0 0 4720 782
4 QDFF
-14 -44 14 -36
3 U16
-57 -4 -36 4
0
15 DVCC=16;DGND=8;
85 %D [%16bi %8bi %1i %2i %3i %4i %9i]
+ [%16bo %1o %2o %3o %4o %9o %5o %6o %7o %8o] %M
0
11 typeDigital
5 DIP16
19

0 1 2 3 4 5 6 7 8 9
1 2 3 4 5 6 7 8 9 0
65 0 0 0 1 0 0 0
1 U
3976 0 0
2
44331.3 72
0
5 7412~
219 1383 878 0 4 22
0 101 399 381 402
0
0 0 624 0
4 7412
-7 -24 21 -16
4 U15A
-15 -12 13 -4
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 3 4 5 6 3 4 5 6 1
2 8 9 11 12 13 10 0 0 0
0 6 0
65 0 0 0 3 1 7 0
1 U
3624 0 0
2
44331.3 73
0
12 D Flip-Flop~
219 1075 338 0 4 9
0 125 124 418 104
0
0 0 4720 0
3 DFF
-10 -53 11 -45
3 U21
-11 -55 10 -47
0
14 DVCC=6;DGND=5;
47 %D [%6bi %5bi %1i %2i][%6bo %1o %2o %3o %4o] %M
0
11 typeDigital
4 DIP6
9

0 1 2 3 4 1 2 3 4 0
65 0 0 512 1 0 0 0
1 U
3912 0 0
2
44331.3 74
0
12 D Flip-Flop~
219 902 331 0 4 9
0 137 136 419 62
0
0 0 4720 0
3 DFF
-10 -53 11 -45
3 U25
-11 -55 10 -47
0
14 DVCC=6;DGND=5;
47 %D [%6bi %5bi %1i %2i][%6bo %1o %2o %3o %4o] %M
0
11 typeDigital
4 DIP6
9

0 1 2 3 4 1 2 3 4 0
65 0 0 512 1 0 0 0
1 U
3928 0 0
2
44331.3 75
0
9 2-In AND~
219 1212 356 0 3 22
0 62 385 103
0
0 0 624 0
6 74LS08
-21 -24 21 -16
4 U12A
-12 -13 16 -5
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 3 0
1 U
4866 0 0
2
44331.3 76
0
6 74266~
219 1130 373 0 3 22
0 104 382 385
0
0 0 624 0
7 74LS266
-24 -24 25 -16
4 U11A
-3 -12 25 -4
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 6 0
1 U
9491 0 0
2
44331.3 77
0
9 Inverter~
13 612 735 0 2 22
0 381 392
0
0 0 624 0
6 74LS04
-21 -19 21 -11
3 U3C
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 5 6 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 3 1 0
1 U
3166 0 0
2
44331.3 78
0
9 Inverter~
13 564 614 0 2 22
0 380 2
0
0 0 624 0
6 74LS04
-21 -19 21 -11
3 U3B
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 3 4 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 2 1 0
1 U
6131 0 0
2
44331.3 79
0
9 Inverter~
13 565 555 0 2 22
0 3 403
0
0 0 624 0
6 74LS04
-21 -19 21 -11
3 U3A
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 1 1 0
1 U
5864 0 0
2
44331.3 80
0
9 2-In AND~
219 663 683 0 3 22
0 3 380 393
0
0 0 624 0
6 74LS08
-21 -24 21 -16
4 U10D
-16 -11 12 -3
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 5 0
1 U
5373 0 0
2
44331.3 81
0
9 2-In AND~
219 663 646 0 3 22
0 3 2 396
0
0 0 624 0
6 74LS08
-21 -24 21 -16
4 U10C
-16 -11 12 -3
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 5 0
1 U
9688 0 0
2
44331.3 82
0
9 2-In AND~
219 663 600 0 3 22
0 403 380 399
0
0 0 624 0
6 74LS08
-21 -24 21 -16
4 U10B
-16 -11 12 -3
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 5 0
1 U
5140 0 0
2
44331.3 83
0
9 2-In AND~
219 663 564 0 3 22
0 403 2 400
0
0 0 624 0
6 74LS08
-21 -24 21 -16
4 U10A
-16 -11 12 -3
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 5 0
1 U
955 0 0
2
44331.3 84
0
5 7412~
219 1375 456 0 4 22
0 103 400 381 404
0
0 0 624 0
4 7412
-7 -24 21 -16
3 U9B
-13 -11 8 -3
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 1 2 8 9 3 4 5 6 1
2 8 9 11 12 13 10 0 0 0
0 6 0
65 0 0 0 3 2 4 0
1 U
3525 0 0
2
44331.3 85
0
5 7412~
219 1289 408 0 4 22
0 103 400 392 405
0
0 0 624 0
4 7412
-7 -24 21 -16
3 U9A
-15 -12 6 -4
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 3 4 5 6 3 4 5 6 1
2 8 9 11 12 13 10 0 0 0
0 6 0
65 0 0 0 3 1 4 0
1 U
4450 0 0
2
44331.3 86
0
12 Quad D Flop~
47 1374 251 0 9 19
0 57 56 55 54 40 39 38 37 161
0
0 0 4720 782
4 QDFF
-14 -44 14 -36
2 U1
-54 -4 -40 4
0
15 DVCC=16;DGND=8;
85 %D [%16bi %8bi %1i %2i %3i %4i %9i]
+ [%16bo %1o %2o %3o %4o %9o %5o %6o %7o %8o] %M
0
11 typeDigital
5 DIP16
19

0 1 2 3 4 5 6 7 8 9
1 2 3 4 5 6 7 8 9 0
65 0 0 0 1 0 0 0
1 U
390 0 0
2
44331.3 87
0
13 Quad 3-State~
48 1377 328 0 9 19
0 40 39 38 37 90 89 88 87 405
0
0 0 4720 782
8 QUAD3STA
-28 -44 28 -36
2 U2
-57 -1 -43 7
0
15 DVCC=16;DGND=8;
85 %D [%16bi %8bi %1i %2i %3i %4i %9i]
+ [%16bo %1o %2o %3o %4o %9o %5o %6o %7o %8o] %M
0
12 type:digital
5 DIP16
19

0 1 2 3 4 5 6 7 8 9
1 2 3 4 5 6 7 8 9 0
65 0 0 0 1 0 0 0
1 U
8631 0 0
2
44331.3 88
0
12 Quad D Flop~
47 1571 256 0 9 19
0 53 52 51 50 24 23 22 21 160
0
0 0 4720 782
4 QDFF
-14 -44 14 -36
2 U7
-54 -4 -40 4
0
15 DVCC=16;DGND=8;
85 %D [%16bi %8bi %1i %2i %3i %4i %9i]
+ [%16bo %1o %2o %3o %4o %9o %5o %6o %7o %8o] %M
0
11 typeDigital
5 DIP16
19

0 1 2 3 4 5 6 7 8 9
1 2 3 4 5 6 7 8 9 0
65 0 0 0 1 0 0 0
1 U
3384 0 0
2
44331.3 89
0
13 Quad 3-State~
48 1574 335 0 9 19
0 24 23 22 21 86 85 84 83 404
0
0 0 4720 782
8 QUAD3STA
-28 -44 28 -36
2 U8
-57 -1 -43 7
0
15 DVCC=16;DGND=8;
85 %D [%16bi %8bi %1i %2i %3i %4i %9i]
+ [%16bo %1o %2o %3o %4o %9o %5o %6o %7o %8o] %M
0
12 type:digital
5 DIP16
19

0 1 2 3 4 5 6 7 8 9
1 2 3 4 5 6 7 8 9 0
65 0 0 0 1 0 0 0
1 U
3527 0 0
2
44331.3 90
0
7 Pulser~
4 645 99 0 10 12
0 420 421 117 422 0 0 5 5 4
7
0
0 0 4656 0
0
2 V5
-7 -28 7 -20
0
0
0
0
0
4 SIP2
9

0 1 2 3 4 1 2 3 4 0
0 0 0 512 1 0 0 0
1 V
3353 0 0
2
44331.3 91
0
642
2 0 2 0 0 8320 0 381 0 0 631 4
639 655
589 655
589 593
585 593
1 0 3 0 0 4096 0 381 0 0 625 2
639 637
533 637
1 0 4 0 0 4096 0 74 0 0 232 2
2869 2547
2869 2496
1 0 5 0 0 4096 0 75 0 0 228 2
2866 2220
2866 2166
1 0 6 0 0 4096 0 76 0 0 224 4
2865 1899
2865 1864
2880 1864
2880 1849
1 0 7 0 0 4096 0 77 0 0 219 2
2874 1594
2874 1543
0 0 8 0 0 12288 0 0 0 112 111 5
2855 629
2837 629
2837 618
2809 618
2809 629
1 0 9 0 0 8320 0 81 0 0 570 3
1756 1593
1756 1624
1590 1624
1 0 10 0 0 8320 0 80 0 0 571 3
1740 1593
1740 1619
1578 1619
1 0 11 0 0 8320 0 79 0 0 572 3
1724 1593
1724 1614
1566 1614
0 1 12 0 0 4224 0 0 78 573 0 3
1554 1609
1708 1609
1708 1593
1 0 13 0 0 8320 0 85 0 0 590 3
1754 1072
1754 1103
1588 1103
1 0 14 0 0 8320 0 84 0 0 591 3
1738 1072
1738 1098
1576 1098
1 0 15 0 0 8320 0 83 0 0 592 3
1722 1072
1722 1093
1564 1093
0 1 16 0 0 4224 0 0 82 593 0 3
1552 1088
1706 1088
1706 1072
1 0 17 0 0 8320 0 89 0 0 611 3
1749 680
1749 711
1583 711
1 0 18 0 0 8320 0 88 0 0 612 3
1733 680
1733 706
1571 706
1 0 19 0 0 8320 0 87 0 0 613 3
1717 680
1717 701
1559 701
0 1 20 0 0 4224 0 0 86 614 0 3
1547 696
1701 696
1701 680
1 0 21 0 0 8320 0 90 0 0 635 3
1743 273
1743 304
1577 304
1 0 22 0 0 8320 0 91 0 0 636 3
1727 273
1727 299
1565 299
1 0 23 0 0 8320 0 92 0 0 637 3
1711 273
1711 294
1553 294
0 1 24 0 0 4224 0 0 93 638 0 3
1541 289
1695 289
1695 273
1 0 25 0 0 8320 0 97 0 0 565 3
1325 1598
1325 1620
1400 1620
1 0 26 0 0 8320 0 96 0 0 566 3
1309 1598
1309 1614
1388 1614
1 0 27 0 0 8320 0 95 0 0 567 3
1293 1598
1293 1609
1376 1609
1 0 28 0 0 8320 0 94 0 0 568 3
1277 1598
1277 1606
1364 1606
1 0 29 0 0 8320 0 101 0 0 585 3
1318 1078
1318 1100
1393 1100
1 0 30 0 0 8320 0 100 0 0 586 3
1302 1078
1302 1094
1381 1094
1 0 31 0 0 8320 0 99 0 0 587 3
1286 1078
1286 1089
1369 1089
1 0 32 0 0 8320 0 98 0 0 588 3
1270 1078
1270 1086
1357 1086
1 0 33 0 0 8320 0 105 0 0 606 3
1309 685
1309 707
1384 707
1 0 34 0 0 8320 0 104 0 0 607 3
1293 685
1293 701
1372 701
1 0 35 0 0 8320 0 103 0 0 608 3
1277 685
1277 696
1360 696
1 0 36 0 0 8320 0 102 0 0 609 3
1261 685
1261 693
1348 693
1 0 37 0 0 8320 0 106 0 0 639 3
1305 274
1305 296
1380 296
1 0 38 0 0 8320 0 107 0 0 640 3
1289 274
1289 290
1368 290
1 0 39 0 0 8320 0 108 0 0 641 3
1273 274
1273 285
1356 285
1 0 40 0 0 8320 0 109 0 0 642 3
1257 274
1257 282
1344 282
5 5 41 0 0 12416 0 337 342 0 0 4
1513 2016
1541 2016
1541 2034
1589 2034
3 1 42 0 0 8320 0 180 110 0 0 3
1687 1827
1640 1827
1640 1769
3 2 43 0 0 4224 0 179 110 0 0 3
1687 1789
1658 1789
1658 1769
0 0 44 0 0 8320 0 0 0 189 120 4
1452 1255
1452 1259
883 1259
883 1146
2 3 45 0 0 4224 0 111 181 0 0 3
1660 1237
1660 1296
1719 1296
3 1 46 0 0 4224 0 182 111 0 0 3
1718 1262
1642 1262
1642 1237
0 0 47 0 0 8320 0 0 0 201 122 4
1436 434
1436 433
846 433
846 357
3 2 48 0 0 4224 0 183 112 0 0 4
1706 868
1656 868
1656 818
1654 818
1 3 49 0 0 8320 0 112 184 0 0 3
1636 818
1636 833
1706 833
4 3 50 0 0 4224 0 388 229 0 0 3
1577 232
1610 232
1610 216
3 3 51 0 0 4224 0 388 228 0 0 3
1565 232
1565 216
1577 216
3 2 52 0 0 8320 0 227 388 0 0 3
1544 216
1553 216
1553 232
3 1 53 0 0 8320 0 230 388 0 0 4
1511 215
1511 224
1541 224
1541 232
4 3 54 0 0 8320 0 386 232 0 0 4
1380 227
1380 225
1413 225
1413 214
3 3 55 0 0 8320 0 233 386 0 0 4
1380 212
1380 219
1368 219
1368 227
3 2 56 0 0 8320 0 329 386 0 0 4
1347 212
1347 219
1356 219
1356 227
3 1 57 0 0 8320 0 231 386 0 0 4
1314 212
1314 219
1344 219
1344 227
2 3 58 0 0 8320 0 114 185 0 0 3
1658 405
1658 453
1712 453
3 1 59 0 0 4224 0 186 114 0 0 3
1712 418
1640 418
1640 405
0 0 60 0 0 4096 0 0 0 114 139 2
2811 332
2850 332
1 0 61 0 0 4096 0 115 0 0 603 2
948 694
948 693
1 0 62 0 0 0 0 116 0 0 622 2
939 295
939 295
8 1 63 0 0 8320 0 352 118 0 0 3
1590 1713
1599 1713
1599 1730
7 1 64 0 0 8320 0 352 117 0 0 3
1578 1713
1583 1713
1583 1730
1 6 65 0 0 12416 0 119 352 0 0 4
1567 1730
1567 1722
1566 1722
1566 1713
5 1 66 0 0 8320 0 352 120 0 0 3
1554 1713
1551 1713
1551 1730
8 1 67 0 0 8320 0 347 122 0 0 3
1400 1713
1409 1713
1409 1730
7 1 68 0 0 8320 0 347 121 0 0 3
1388 1713
1393 1713
1393 1730
1 6 69 0 0 4224 0 123 347 0 0 3
1377 1730
1377 1713
1376 1713
5 1 70 0 0 8320 0 347 124 0 0 3
1364 1713
1361 1713
1361 1730
8 1 71 0 0 8320 0 362 126 0 0 3
1588 1183
1597 1183
1597 1197
7 1 72 0 0 8320 0 362 125 0 0 3
1576 1183
1581 1183
1581 1197
1 6 73 0 0 4224 0 127 362 0 0 3
1565 1197
1565 1183
1564 1183
5 1 74 0 0 8320 0 362 128 0 0 3
1552 1183
1549 1183
1549 1197
8 1 75 0 0 8320 0 357 130 0 0 3
1393 1181
1402 1181
1402 1198
7 1 76 0 0 8320 0 357 129 0 0 3
1381 1181
1386 1181
1386 1198
1 6 77 0 0 12416 0 131 357 0 0 4
1370 1198
1370 1190
1369 1190
1369 1181
5 1 78 0 0 8320 0 357 132 0 0 3
1357 1181
1354 1181
1354 1198
8 1 79 0 0 8320 0 370 134 0 0 3
1583 775
1592 775
1592 786
7 1 80 0 0 8320 0 370 133 0 0 3
1571 775
1576 775
1576 786
1 6 81 0 0 4224 0 135 370 0 0 3
1560 786
1560 775
1559 775
5 1 82 0 0 8320 0 370 136 0 0 3
1547 775
1544 775
1544 786
8 1 83 0 0 4224 0 389 138 0 0 3
1577 362
1586 362
1586 368
7 1 84 0 0 8320 0 389 137 0 0 3
1565 362
1570 362
1570 368
1 6 85 0 0 4224 0 139 389 0 0 4
1554 368
1554 365
1553 365
1553 362
5 1 86 0 0 8320 0 389 140 0 0 3
1541 362
1538 362
1538 368
8 1 87 0 0 8320 0 387 142 0 0 3
1380 355
1389 355
1389 366
7 1 88 0 0 8320 0 387 141 0 0 3
1368 355
1373 355
1373 366
1 6 89 0 0 12416 0 143 387 0 0 4
1357 366
1357 361
1356 361
1356 355
5 1 90 0 0 8320 0 387 144 0 0 3
1344 355
1341 355
1341 366
8 1 91 0 0 8320 0 369 147 0 0 3
1384 774
1394 774
1394 788
7 1 92 0 0 8320 0 369 148 0 0 3
1372 774
1378 774
1378 788
1 6 93 0 0 4224 0 146 369 0 0 4
1363 788
1363 781
1360 781
1360 774
5 1 94 0 0 4224 0 369 145 0 0 2
1348 774
1348 788
1 0 95 0 0 0 0 149 0 0 527 2
1294 1695
1294 1695
1 0 96 0 0 4096 0 150 0 0 562 2
1142 1603
1145 1603
1 0 97 0 0 4096 0 151 0 0 563 2
986 1606
989 1606
1 0 98 0 0 0 0 152 0 0 580 2
1278 1140
1278 1140
1 0 99 0 0 4096 0 153 0 0 582 2
967 1068
967 1070
1 0 100 0 0 0 0 154 0 0 581 2
1144 1073
1144 1073
1 0 101 0 0 0 0 155 0 0 601 2
1256 758
1256 758
1 0 102 0 0 0 0 156 0 0 602 2
1120 696
1120 696
1 0 103 0 0 4096 0 157 0 0 621 2
1257 356
1258 356
1 0 104 0 0 4096 0 158 0 0 620 2
1111 302
1112 302
2 0 105 0 0 8320 0 159 0 0 0 5
1029 1505
1029 1366
2323 1366
2323 1276
2822 1276
2 1 106 0 0 8320 0 74 159 0 0 5
2833 2547
1940 2547
1940 1381
1047 1381
1047 1505
1 2 107 0 0 12416 0 160 75 0 0 5
1035 972
1035 939
2246 939
2246 2220
2830 2220
0 2 108 0 0 12416 0 0 160 0 0 5
2840 939
2276 939
2276 929
1017 929
1017 972
2 1 109 0 0 8320 0 76 161 0 0 5
2829 1899
2091 1899
2091 522
1017 522
1017 581
0 0 105 0 0 0 0 0 0 104 217 6
2807 1276
2807 1269
2841 1269
2841 1276
2862 1276
2862 1226
0 0 108 0 0 0 0 0 0 107 213 6
2830 939
2830 926
2867 926
2867 939
2880 939
2880 889
0 2 8 0 0 4224 0 0 161 0 0 5
2816 629
1904 629
1904 492
999 492
999 581
0 0 8 0 0 0 0 0 0 212 0 3
2855 582
2855 629
2852 629
2 1 110 0 0 8320 0 77 162 0 0 5
2838 1594
2086 1594
2086 74
1014 74
1014 186
2 0 60 0 0 8320 0 162 0 0 0 4
996 186
996 64
2811 64
2811 341
1 3 111 0 0 8320 0 164 159 0 0 4
1022 1584
1009 1584
1009 1551
1038 1551
3 1 112 0 0 8320 0 160 166 0 0 4
1026 1018
1001 1018
1001 1054
1022 1054
1 3 113 0 0 8320 0 168 161 0 0 5
998 677
977 677
977 635
1008 635
1008 627
1 3 114 0 0 8320 0 169 162 0 0 5
988 283
979 283
979 244
1005 244
1005 232
0 0 115 0 0 8192 0 0 0 126 145 3
1043 1645
1043 1679
894 1679
0 0 44 0 0 0 0 0 0 129 150 4
1044 1115
1044 1146
882 1146
882 1108
0 0 116 0 0 8192 0 0 0 132 154 3
1020 738
1020 771
860 771
0 0 47 0 0 0 0 0 0 159 136 4
846 333
846 360
1008 360
1008 342
1 0 117 0 0 8192 0 163 0 0 124 3
1008 1629
997 1629
997 1099
1 0 117 0 0 0 0 165 0 0 125 5
1008 1099
977 1099
977 759
968 759
968 722
1 0 117 0 0 0 0 167 0 0 135 3
984 722
961 722
961 328
2 2 115 0 0 0 0 164 163 0 0 5
1037 1595
1054 1595
1054 1645
1023 1645
1023 1640
3 2 118 0 0 4224 0 163 343 0 0 4
1038 1629
1071 1629
1071 1621
1084 1621
3 1 119 0 0 8320 0 164 343 0 0 4
1052 1584
1070 1584
1070 1603
1084 1603
2 2 44 0 0 0 0 166 165 0 0 5
1037 1065
1054 1065
1054 1115
1023 1115
1023 1110
3 2 120 0 0 4224 0 165 353 0 0 4
1038 1099
1071 1099
1071 1091
1084 1091
3 1 121 0 0 8320 0 166 353 0 0 4
1052 1054
1070 1054
1070 1073
1084 1073
2 2 116 0 0 0 0 168 167 0 0 5
1013 688
1030 688
1030 738
999 738
999 733
3 2 122 0 0 4224 0 167 366 0 0 4
1014 722
1047 722
1047 714
1060 714
3 1 123 0 0 8320 0 168 366 0 0 4
1028 677
1046 677
1046 696
1060 696
1 0 117 0 0 0 0 170 0 0 199 3
974 328
952 328
952 90
2 2 47 0 0 0 0 169 170 0 0 5
1003 294
1020 294
1020 342
989 342
989 339
3 2 124 0 0 4224 0 170 373 0 0 4
1004 328
1037 328
1037 320
1051 320
3 1 125 0 0 8320 0 169 373 0 0 4
1018 283
1036 283
1036 302
1051 302
0 0 60 0 0 0 0 0 0 211 0 3
2850 295
2850 341
2847 341
0 1 117 0 0 4224 0 0 171 141 0 3
772 1095
772 1632
862 1632
0 1 117 0 0 0 0 0 173 142 0 3
772 719
772 1096
850 1096
0 1 117 0 0 0 0 0 175 143 0 3
772 321
772 719
828 719
3 1 117 0 0 0 0 390 178 0 0 4
669 90
771 90
771 321
814 321
1 1 126 0 0 4224 0 1 172 0 0 2
854 1587
862 1587
0 0 115 0 0 8320 0 0 0 187 146 6
1461 1796
1461 1798
1072 1798
1072 1720
894 1720
894 1648
2 2 115 0 0 0 0 172 171 0 0 5
877 1598
894 1598
894 1648
877 1648
877 1643
3 2 127 0 0 4224 0 171 344 0 0 4
892 1632
911 1632
911 1624
925 1624
3 1 128 0 0 8320 0 172 344 0 0 4
892 1587
910 1587
910 1606
925 1606
1 1 129 0 0 4224 0 2 174 0 0 2
842 1051
850 1051
2 2 44 0 0 0 0 174 173 0 0 5
865 1062
882 1062
882 1112
865 1112
865 1107
3 2 130 0 0 4224 0 173 354 0 0 4
880 1096
899 1096
899 1088
913 1088
3 1 131 0 0 8320 0 174 354 0 0 4
880 1051
898 1051
898 1070
913 1070
1 1 132 0 0 4224 0 3 176 0 0 2
820 674
828 674
0 0 116 0 0 8320 0 0 0 195 155 6
1459 856
1459 858
1106 858
1106 816
860 816
860 735
2 2 116 0 0 0 0 176 175 0 0 5
843 685
860 685
860 735
843 735
843 730
3 2 133 0 0 4224 0 175 365 0 0 4
858 719
877 719
877 711
891 711
3 1 134 0 0 8320 0 176 365 0 0 4
858 674
876 674
876 693
891 693
1 1 135 0 0 4224 0 4 177 0 0 2
806 276
814 276
2 2 47 0 0 0 0 177 178 0 0 5
829 287
846 287
846 337
829 337
829 332
3 2 136 0 0 4224 0 178 374 0 0 4
844 321
863 321
863 313
878 313
3 1 137 0 0 8320 0 177 374 0 0 4
844 276
862 276
862 295
878 295
22 1 138 0 0 8192 0 342 180 0 0 4
1653 2106
1815 2106
1815 1836
1733 1836
0 1 139 0 0 8192 0 0 179 230 0 4
1665 2097
1820 2097
1820 1798
1733 1798
1 0 140 0 0 8192 0 181 0 0 227 4
1765 1305
2117 1305
2117 2088
1675 2088
0 1 141 0 0 8192 0 0 182 226 0 4
1685 2079
2125 2079
2125 1271
1764 1271
1 0 142 0 0 8192 0 183 0 0 223 4
1752 877
2133 877
2133 2070
1691 2070
0 1 143 0 0 8192 0 0 184 222 0 4
1702 2061
2137 2061
2137 842
1752 842
1 0 144 0 0 8320 0 185 0 0 221 4
1758 462
2142 462
2142 2052
1711 2052
1 0 145 0 0 8320 0 186 0 0 210 4
1758 427
2148 427
2148 2043
1724 2043
0 2 146 0 0 8192 0 0 180 209 0 4
1734 2034
1826 2034
1826 1818
1733 1818
0 2 147 0 0 8192 0 0 179 208 0 4
1743 2025
1834 2025
1834 1780
1733 1780
0 1 117 0 0 0 0 0 187 182 0 3
1682 1054
1682 1574
1658 1574
0 1 117 0 0 0 0 0 188 183 0 4
1490 1054
1480 1054
1480 1570
1470 1570
3 9 148 0 0 4224 0 187 351 0 0 4
1628 1574
1624 1574
1624 1573
1620 1573
3 9 149 0 0 4224 0 188 348 0 0 2
1440 1570
1430 1570
0 2 150 0 0 8192 0 0 181 207 0 4
1753 2016
2234 2016
2234 1287
1765 1287
0 2 151 0 0 8192 0 0 182 206 0 4
1762 2007
2222 2007
2222 1253
1764 1253
2 0 152 0 0 4096 0 183 0 0 205 2
1752 859
2213 859
2 0 153 0 0 4096 0 184 0 0 204 2
1752 824
2203 824
2 0 154 0 0 4096 0 185 0 0 203 2
1758 444
2195 444
2 0 155 0 0 4096 0 186 0 0 202 2
1758 409
2188 409
0 1 117 0 0 0 0 0 189 190 0 3
1682 661
1682 1056
1656 1056
1 0 117 0 0 0 0 190 0 0 192 4
1459 1054
1490 1054
1490 662
1470 662
3 9 156 0 0 4224 0 189 361 0 0 2
1626 1056
1618 1056
3 9 157 0 0 4224 0 190 358 0 0 4
1429 1054
1425 1054
1425 1050
1423 1050
3 2 115 0 0 0 0 110 187 0 0 4
1649 1723
1649 1598
1643 1598
1643 1585
0 2 115 0 0 0 0 0 188 186 0 7
1649 1696
1631 1696
1631 1796
1458 1796
1458 1599
1455 1599
1455 1581
3 2 44 0 0 0 0 111 189 0 0 4
1651 1191
1651 1075
1641 1075
1641 1067
0 2 44 0 0 0 0 0 190 188 0 7
1651 1170
1631 1170
1631 1255
1452 1255
1452 1076
1444 1076
1444 1065
0 1 117 0 0 0 0 0 191 196 0 4
1647 243
1682 243
1682 661
1660 661
3 9 158 0 0 4224 0 191 371 0 0 2
1630 661
1613 661
1 0 117 0 0 0 0 192 0 0 199 4
1447 662
1472 662
1472 237
1456 237
3 9 159 0 0 4224 0 192 368 0 0 2
1417 662
1414 662
3 2 116 0 0 0 0 112 191 0 0 2
1645 772
1645 672
0 2 116 0 0 0 0 0 192 194 0 7
1645 761
1624 761
1624 856
1458 856
1458 686
1432 686
1432 673
0 1 117 0 0 0 0 0 193 199 0 4
1456 91
1647 91
1647 256
1642 256
3 9 160 0 0 4224 0 193 388 0 0 2
1612 256
1607 256
3 2 47 0 0 0 0 114 193 0 0 4
1649 359
1649 284
1627 284
1627 267
1 0 117 0 0 0 0 194 0 0 143 7
1444 251
1444 237
1456 237
1456 89
1061 89
1061 90
771 90
3 9 161 0 0 4224 0 194 386 0 0 2
1414 251
1410 251
0 2 47 0 0 0 0 0 194 198 0 7
1649 344
1625 344
1625 434
1436 434
1436 283
1429 283
1429 262
7 2 155 0 0 8320 0 342 202 0 0 6
1653 1971
2188 1971
2188 361
2944 361
2944 286
2931 286
8 1 154 0 0 8320 0 342 202 0 0 6
1653 1980
2195 1980
2195 367
2938 367
2938 304
2931 304
9 2 153 0 0 8320 0 342 201 0 0 6
1653 1989
2203 1989
2203 653
2957 653
2957 573
2929 573
10 1 152 0 0 8320 0 342 201 0 0 6
1653 1998
2213 1998
2213 644
2942 644
2942 591
2929 591
11 2 151 0 0 16512 0 342 200 0 0 6
1653 2007
1762 2007
1762 2627
3022 2627
3022 880
2938 880
12 1 150 0 0 16512 0 342 200 0 0 6
1653 2016
1753 2016
1753 2631
3019 2631
3019 898
2938 898
13 2 147 0 0 16512 0 342 199 0 0 6
1653 2025
1743 2025
1743 2635
3013 2635
3013 1217
2917 1217
14 1 146 0 0 16512 0 342 199 0 0 6
1653 2034
1734 2034
1734 2639
3008 2639
3008 1235
2917 1235
15 2 145 0 0 0 0 342 198 0 0 6
1653 2043
1724 2043
1724 2641
3005 2641
3005 1534
2943 1534
3 0 60 0 0 0 0 202 0 0 216 2
2879 295
2777 295
3 0 8 0 0 0 0 201 0 0 215 2
2877 582
2780 582
3 0 108 0 0 0 0 200 0 0 214 2
2886 889
2784 889
9 9 108 0 0 0 0 308 317 0 0 4
2497 850
2497 910
2784 910
2784 842
9 9 8 0 0 0 0 256 247 0 0 4
2493 548
2493 603
2780 603
2780 540
9 9 60 0 0 0 0 330 320 0 0 4
2490 267
2490 319
2777 319
2777 259
3 0 105 0 0 0 0 199 0 0 218 2
2865 1226
2785 1226
9 9 105 0 0 0 0 296 305 0 0 4
2498 1186
2498 1235
2785 1235
2785 1178
3 0 7 0 0 4096 0 198 0 0 220 2
2891 1543
2791 1543
9 9 7 0 0 8320 0 244 235 0 0 4
2504 1495
2504 1606
2791 1606
2791 1487
16 1 144 0 0 0 0 342 198 0 0 6
1653 2052
1713 2052
1713 2643
3002 2643
3002 1552
2943 1552
17 2 143 0 0 12416 0 342 197 0 0 6
1653 2061
1703 2061
1703 2647
2996 2647
2996 1840
2944 1840
18 1 142 0 0 12416 0 342 197 0 0 6
1653 2070
1693 2070
1693 2649
2991 2649
2991 1858
2944 1858
3 0 6 0 0 4096 0 197 0 0 225 2
2892 1849
2795 1849
9 9 6 0 0 12416 0 269 260 0 0 5
2508 1808
2556 1808
2556 1914
2795 1914
2795 1800
19 2 141 0 0 12416 0 342 196 0 0 6
1653 2079
1685 2079
1685 2653
2988 2653
2988 2157
2946 2157
20 1 140 0 0 12416 0 342 196 0 0 6
1653 2088
1675 2088
1675 2656
2981 2656
2981 2175
2946 2175
3 0 5 0 0 4096 0 196 0 0 229 2
2894 2166
2792 2166
9 9 5 0 0 12416 0 281 272 0 0 5
2505 2124
2550 2124
2550 2235
2792 2235
2792 2116
21 2 139 0 0 12416 0 342 195 0 0 6
1653 2097
1665 2097
1665 2661
2974 2661
2974 2487
2946 2487
22 1 138 0 0 8320 0 342 195 0 0 5
1653 2106
1653 2668
2969 2668
2969 2505
2946 2505
3 0 4 0 0 4096 0 195 0 0 233 2
2894 2496
2793 2496
9 9 4 0 0 12416 0 293 284 0 0 5
2506 2460
2551 2460
2551 2564
2793 2564
2793 2452
0 9 162 0 0 4224 0 0 283 236 0 3
2807 2057
2807 2395
2787 2395
9 0 162 0 0 0 0 294 0 0 237 3
2500 2403
2534 2403
2534 2067
0 9 162 0 0 0 0 0 271 238 0 3
2807 1743
2807 2059
2786 2059
9 0 162 0 0 0 0 282 0 0 239 4
2499 2067
2534 2067
2534 1743
2517 1743
9 0 162 0 0 0 0 259 0 0 240 4
2789 1743
2808 1743
2808 1430
2794 1430
0 9 162 0 0 0 0 0 270 241 0 4
2524 1433
2517 1433
2517 1751
2502 1751
0 9 162 0 0 0 0 0 234 242 0 3
2794 1121
2794 1430
2785 1430
0 9 162 0 0 0 0 0 245 243 0 4
2520 1129
2524 1129
2524 1438
2498 1438
9 0 162 0 0 0 0 306 0 0 244 3
2779 1121
2794 1121
2794 783
0 9 162 0 0 0 0 0 295 245 0 4
2518 793
2520 793
2520 1129
2492 1129
0 9 162 0 0 0 0 0 318 246 0 3
2794 483
2794 785
2778 785
9 0 162 0 0 0 0 307 0 0 247 4
2491 793
2518 793
2518 487
2505 487
9 0 162 0 0 0 0 246 0 0 249 3
2774 483
2794 483
2794 202
9 0 162 0 0 0 0 257 0 0 249 3
2487 491
2505 491
2505 205
3 0 162 0 0 0 0 258 0 0 249 4
2895 33
2930 33
2930 72
2794 72
9 9 162 0 0 0 0 331 319 0 0 6
2484 210
2505 210
2505 72
2794 72
2794 202
2771 202
1 8 163 0 0 12416 0 204 284 0 0 6
1632 1485
1632 1470
1841 1470
1841 2532
2757 2532
2757 2476
7 1 164 0 0 12416 0 284 205 0 0 6
2745 2476
2745 2527
1849 2527
1849 1466
1599 1466
1599 1485
1 6 165 0 0 12416 0 206 284 0 0 6
1566 1484
1566 1456
1856 1456
1856 2518
2733 2518
2733 2476
5 1 166 0 0 12416 0 284 203 0 0 6
2721 2476
2721 2515
1861 2515
1861 1449
1533 1449
1533 1484
1 8 167 0 0 12416 0 208 293 0 0 6
1442 1482
1442 1444
1870 1444
1870 2509
2470 2509
2470 2484
7 1 168 0 0 12416 0 293 209 0 0 6
2458 2484
2458 2501
1874 2501
1874 1436
1409 1436
1409 1482
1 6 169 0 0 12416 0 210 293 0 0 6
1376 1481
1376 1429
1879 1429
1879 2493
2446 2493
2446 2484
5 1 170 0 0 8320 0 293 207 0 0 5
2434 2484
1883 2484
1883 1421
1343 1421
1343 1481
1 8 171 0 0 8320 0 212 272 0 0 5
1630 968
1893 968
1893 2206
2756 2206
2756 2140
7 1 172 0 0 12416 0 272 213 0 0 6
2744 2140
2744 2199
1901 2199
1901 961
1597 961
1597 968
6 1 173 0 0 12416 0 272 214 0 0 6
2732 2140
2732 2194
1907 2194
1907 956
1564 956
1564 967
5 1 174 0 0 12416 0 272 211 0 0 6
2720 2140
2720 2191
1911 2191
1911 952
1531 952
1531 967
8 1 175 0 0 12416 0 281 216 0 0 6
2469 2148
2469 2166
1917 2166
1917 948
1435 948
1435 966
1 7 176 0 0 12416 0 217 281 0 0 6
1402 966
1402 942
1919 942
1919 2161
2457 2161
2457 2148
6 1 177 0 0 12416 0 281 218 0 0 6
2445 2148
2445 2154
1922 2154
1922 936
1369 936
1369 965
5 1 178 0 0 8320 0 281 215 0 0 5
2433 2148
1925 2148
1925 932
1336 932
1336 965
1 8 179 0 0 12416 0 220 260 0 0 6
1625 573
1625 560
1955 560
1955 1894
2759 1894
2759 1824
7 1 180 0 0 12416 0 260 221 0 0 6
2747 1824
2747 1886
1961 1886
1961 555
1592 555
1592 573
6 1 181 0 0 12416 0 260 222 0 0 6
2735 1824
2735 1876
1967 1876
1967 549
1559 549
1559 572
5 1 182 0 0 12416 0 260 219 0 0 6
2723 1824
2723 1868
1972 1868
1972 541
1526 541
1526 572
1 8 183 0 0 12416 0 224 269 0 0 6
1426 574
1426 532
1991 532
1991 1856
2472 1856
2472 1832
7 1 184 0 0 12416 0 269 225 0 0 6
2460 1832
2460 1850
2000 1850
2000 525
1393 525
1393 574
6 1 185 0 0 12416 0 269 226 0 0 6
2448 1832
2448 1844
2005 1844
2005 518
1360 518
1360 573
5 1 186 0 0 12416 0 269 223 0 0 6
2436 1832
2436 1841
2012 1841
2012 514
1327 514
1327 573
8 1 187 0 0 12416 0 235 229 0 0 6
2755 1511
2755 1589
2044 1589
2044 164
1619 164
1619 170
7 1 188 0 0 12416 0 235 228 0 0 6
2743 1511
2743 1582
2048 1582
2048 155
1586 155
1586 170
6 1 189 0 0 12416 0 235 227 0 0 6
2731 1511
2731 1573
2052 1573
2052 146
1553 146
1553 170
5 1 190 0 0 12416 0 235 230 0 0 6
2719 1511
2719 1565
2057 1565
2057 136
1520 136
1520 169
1 8 191 0 0 12416 0 232 244 0 0 6
1422 168
1422 130
2072 130
2072 1556
2468 1556
2468 1519
7 1 192 0 0 12416 0 244 233 0 0 6
2456 1519
2456 1546
2074 1546
2074 123
1389 123
1389 166
6 1 193 0 0 12416 0 244 329 0 0 6
2444 1519
2444 1534
2077 1534
2077 119
1356 119
1356 166
1 5 194 0 0 12416 0 231 244 0 0 6
1323 166
1323 112
2081 112
2081 1523
2432 1523
2432 1519
2 8 195 0 0 16512 0 204 305 0 0 6
1614 1485
1614 1413
1899 1413
1899 1273
2749 1273
2749 1202
2 7 196 0 0 16512 0 205 305 0 0 6
1581 1485
1581 1406
1888 1406
1888 1262
2737 1262
2737 1202
2 6 197 0 0 16512 0 206 305 0 0 6
1548 1484
1548 1399
1876 1399
1876 1254
2725 1254
2725 1202
2 5 198 0 0 16512 0 203 305 0 0 6
1515 1484
1515 1393
1866 1393
1866 1245
2713 1245
2713 1202
2 8 199 0 0 16512 0 208 296 0 0 6
1424 1482
1424 1356
1682 1356
1682 1241
2462 1241
2462 1210
2 7 200 0 0 16512 0 209 296 0 0 6
1391 1482
1391 1345
1862 1345
1862 1236
2450 1236
2450 1210
2 6 201 0 0 16512 0 210 296 0 0 6
1358 1481
1358 1335
1857 1335
1857 1230
2438 1230
2438 1210
2 5 202 0 0 16512 0 207 296 0 0 6
1325 1481
1325 1324
1852 1324
1852 1225
2426 1225
2426 1210
8 4 203 0 0 4224 0 295 296 0 0 2
2462 1153
2462 1162
7 3 204 0 0 4224 0 295 296 0 0 2
2450 1153
2450 1162
6 2 205 0 0 4224 0 295 296 0 0 2
2438 1153
2438 1162
5 1 206 0 0 4224 0 295 296 0 0 2
2426 1153
2426 1162
2 8 207 0 0 8320 0 212 317 0 0 4
1612 968
1612 926
2748 926
2748 866
2 7 208 0 0 8320 0 213 317 0 0 4
1579 968
1579 923
2736 923
2736 866
2 6 209 0 0 8320 0 214 317 0 0 4
1546 967
1546 920
2724 920
2724 866
2 5 210 0 0 8320 0 211 317 0 0 4
1513 967
1513 918
2712 918
2712 866
2 8 211 0 0 8320 0 216 308 0 0 6
1417 966
1417 911
2260 911
2260 894
2461 894
2461 874
2 7 212 0 0 8320 0 217 308 0 0 6
1384 966
1384 906
2250 906
2250 885
2449 885
2449 874
2 6 213 0 0 8320 0 218 308 0 0 6
1351 965
1351 902
2242 902
2242 878
2437 878
2437 874
5 2 214 0 0 12416 0 308 215 0 0 5
2425 874
2237 874
2237 898
1318 898
1318 965
2 8 215 0 0 8320 0 220 247 0 0 6
1607 573
1607 509
2245 509
2245 638
2744 638
2744 564
2 7 216 0 0 8320 0 221 247 0 0 6
1574 573
1574 503
2253 503
2253 632
2732 632
2732 564
2 6 217 0 0 8320 0 222 247 0 0 6
1541 572
1541 500
2260 500
2260 623
2720 623
2720 564
2 5 218 0 0 8320 0 219 247 0 0 6
1508 572
1508 495
2266 495
2266 613
2708 613
2708 564
2 8 219 0 0 8320 0 224 256 0 0 6
1408 574
1408 489
2269 489
2269 603
2457 603
2457 572
2 7 220 0 0 8320 0 225 256 0 0 6
1375 574
1375 486
2272 486
2272 598
2445 598
2445 572
2 6 221 0 0 8320 0 226 256 0 0 6
1342 573
1342 481
2275 481
2275 595
2433 595
2433 572
5 2 222 0 0 16512 0 256 223 0 0 6
2421 572
2421 590
2277 590
2277 477
1309 477
1309 573
2 8 223 0 0 8320 0 229 320 0 0 6
1601 170
1601 160
2266 160
2266 357
2741 357
2741 283
2 7 224 0 0 8320 0 228 320 0 0 6
1568 170
1568 151
2273 151
2273 352
2729 352
2729 283
6 2 225 0 0 16512 0 320 227 0 0 6
2717 283
2717 348
2279 348
2279 141
1535 141
1535 170
2 5 226 0 0 8320 0 230 320 0 0 6
1502 169
1502 133
2286 133
2286 344
2705 344
2705 283
2 8 227 0 0 8320 0 232 330 0 0 6
1404 168
1404 126
2290 126
2290 319
2454 319
2454 291
2 7 228 0 0 8320 0 233 330 0 0 6
1371 166
1371 121
2296 121
2296 313
2442 313
2442 291
2 6 229 0 0 8320 0 329 330 0 0 6
1338 166
1338 116
2301 116
2301 305
2430 305
2430 291
2 5 230 0 0 8320 0 231 330 0 0 6
1305 166
1305 109
2305 109
2305 295
2418 295
2418 291
3 3 231 0 0 8320 0 351 205 0 0 4
1578 1549
1578 1538
1590 1538
1590 1531
4 3 232 0 0 8320 0 351 204 0 0 4
1590 1549
1590 1546
1623 1546
1623 1531
3 2 233 0 0 4224 0 206 351 0 0 4
1557 1530
1557 1542
1566 1542
1566 1549
1 3 234 0 0 16512 0 351 203 0 0 6
1554 1549
1554 1545
1543 1545
1543 1531
1524 1531
1524 1530
3 3 235 0 0 8320 0 348 209 0 0 4
1388 1546
1388 1535
1400 1535
1400 1528
4 3 236 0 0 8320 0 348 208 0 0 4
1400 1546
1400 1543
1433 1543
1433 1528
3 2 237 0 0 4224 0 210 348 0 0 4
1367 1527
1367 1539
1376 1539
1376 1546
1 3 238 0 0 16512 0 348 207 0 0 6
1364 1546
1364 1542
1353 1542
1353 1528
1334 1528
1334 1527
3 3 239 0 0 8320 0 361 213 0 0 4
1576 1032
1576 1021
1588 1021
1588 1014
4 3 240 0 0 8320 0 361 212 0 0 4
1588 1032
1588 1029
1621 1029
1621 1014
3 2 241 0 0 4224 0 214 361 0 0 4
1555 1013
1555 1025
1564 1025
1564 1032
1 3 242 0 0 16512 0 361 211 0 0 6
1552 1032
1552 1028
1541 1028
1541 1014
1522 1014
1522 1013
3 3 243 0 0 8320 0 358 217 0 0 4
1381 1026
1381 1019
1393 1019
1393 1012
4 3 244 0 0 8320 0 358 216 0 0 4
1393 1026
1393 1024
1426 1024
1426 1012
3 2 245 0 0 8320 0 218 358 0 0 5
1360 1011
1363 1011
1363 1023
1369 1023
1369 1026
1 3 246 0 0 12416 0 358 215 0 0 5
1357 1026
1346 1026
1346 1012
1327 1012
1327 1011
3 3 247 0 0 8320 0 371 221 0 0 4
1571 637
1571 626
1583 626
1583 619
4 3 248 0 0 8320 0 371 220 0 0 4
1583 637
1583 634
1616 634
1616 619
3 2 249 0 0 4224 0 222 371 0 0 4
1550 618
1550 630
1559 630
1559 637
1 3 250 0 0 16512 0 371 219 0 0 6
1547 637
1547 633
1536 633
1536 619
1517 619
1517 618
3 3 251 0 0 8320 0 368 225 0 0 4
1372 638
1372 627
1384 627
1384 620
4 3 252 0 0 8320 0 368 224 0 0 4
1384 638
1384 635
1417 635
1417 620
3 2 253 0 0 4224 0 226 368 0 0 4
1351 619
1351 631
1360 631
1360 638
1 3 254 0 0 16512 0 368 223 0 0 6
1348 638
1348 634
1337 634
1337 620
1318 620
1318 619
0 1 255 0 0 8320 0 0 234 349 0 3
2664 1379
2664 1406
2719 1406
0 2 256 0 0 8320 0 0 234 348 0 4
2703 1379
2703 1394
2731 1394
2731 1406
0 3 257 0 0 12416 0 0 234 347 0 4
2735 1379
2735 1388
2743 1388
2743 1406
4 0 258 0 0 12416 0 234 0 0 346 4
2755 1406
2755 1397
2767 1397
2767 1379
1 1 258 0 0 0 0 236 5 0 0 4
2758 1378
2767 1378
2767 1379
2774 1379
1 1 257 0 0 0 0 237 6 0 0 2
2725 1379
2741 1379
1 1 256 0 0 0 0 238 7 0 0 2
2694 1379
2710 1379
1 1 255 0 0 0 0 239 8 0 0 2
2659 1379
2675 1379
8 4 259 0 0 4224 0 234 235 0 0 2
2755 1454
2755 1463
7 3 260 0 0 4224 0 234 235 0 0 2
2743 1454
2743 1463
6 2 261 0 0 4224 0 234 235 0 0 2
2731 1454
2731 1463
5 1 262 0 0 4224 0 234 235 0 0 2
2719 1454
2719 1463
0 1 263 0 0 8320 0 0 245 361 0 3
2377 1387
2377 1414
2432 1414
0 2 264 0 0 8320 0 0 245 360 0 4
2416 1387
2416 1402
2444 1402
2444 1414
0 3 265 0 0 12416 0 0 245 359 0 4
2448 1387
2448 1396
2456 1396
2456 1414
4 0 266 0 0 12416 0 245 0 0 358 4
2468 1414
2468 1405
2480 1405
2480 1387
1 1 266 0 0 0 0 243 12 0 0 4
2471 1386
2480 1386
2480 1387
2487 1387
1 1 265 0 0 0 0 242 11 0 0 2
2438 1387
2454 1387
1 1 264 0 0 0 0 241 10 0 0 2
2407 1387
2423 1387
1 1 263 0 0 0 0 240 9 0 0 2
2372 1387
2388 1387
8 4 267 0 0 4224 0 245 244 0 0 2
2468 1462
2468 1471
7 3 268 0 0 4224 0 245 244 0 0 2
2456 1462
2456 1471
6 2 269 0 0 4224 0 245 244 0 0 2
2444 1462
2444 1471
5 1 270 0 0 4224 0 245 244 0 0 2
2432 1462
2432 1471
0 1 271 0 0 8320 0 0 246 373 0 3
2653 432
2653 459
2708 459
0 2 272 0 0 8320 0 0 246 372 0 4
2692 432
2692 447
2720 447
2720 459
0 3 273 0 0 12416 0 0 246 371 0 4
2724 432
2724 441
2732 441
2732 459
4 0 274 0 0 12416 0 246 0 0 370 4
2744 459
2744 450
2756 450
2756 432
1 1 274 0 0 0 0 248 13 0 0 4
2747 431
2756 431
2756 432
2763 432
1 1 273 0 0 0 0 249 14 0 0 2
2714 432
2730 432
1 1 272 0 0 0 0 250 15 0 0 2
2683 432
2699 432
1 1 271 0 0 0 0 251 16 0 0 2
2648 432
2664 432
8 4 275 0 0 4224 0 246 247 0 0 2
2744 507
2744 516
7 3 276 0 0 4224 0 246 247 0 0 2
2732 507
2732 516
6 2 277 0 0 4224 0 246 247 0 0 2
2720 507
2720 516
5 1 278 0 0 4224 0 246 247 0 0 2
2708 507
2708 516
0 1 279 0 0 8320 0 0 257 385 0 3
2366 440
2366 467
2421 467
0 2 280 0 0 8320 0 0 257 384 0 4
2405 440
2405 455
2433 455
2433 467
0 3 281 0 0 12416 0 0 257 383 0 4
2437 440
2437 449
2445 449
2445 467
4 0 282 0 0 12416 0 257 0 0 382 4
2457 467
2457 458
2469 458
2469 440
1 1 282 0 0 0 0 255 20 0 0 4
2460 439
2469 439
2469 440
2476 440
1 1 281 0 0 0 0 254 19 0 0 2
2427 440
2443 440
1 1 280 0 0 0 0 253 18 0 0 2
2396 440
2412 440
1 1 279 0 0 0 0 252 17 0 0 2
2361 440
2377 440
8 4 283 0 0 4224 0 257 256 0 0 2
2457 515
2457 524
7 3 284 0 0 4224 0 257 256 0 0 2
2445 515
2445 524
6 2 285 0 0 4224 0 257 256 0 0 2
2433 515
2433 524
5 1 286 0 0 4224 0 257 256 0 0 2
2421 515
2421 524
0 1 287 0 0 8320 0 0 283 397 0 3
2666 2344
2666 2371
2721 2371
0 2 288 0 0 8320 0 0 283 396 0 4
2705 2344
2705 2359
2733 2359
2733 2371
0 3 289 0 0 12416 0 0 283 395 0 4
2737 2344
2737 2353
2745 2353
2745 2371
4 0 290 0 0 12416 0 283 0 0 394 4
2757 2371
2757 2362
2769 2362
2769 2344
1 1 290 0 0 0 0 285 37 0 0 4
2760 2343
2769 2343
2769 2344
2776 2344
1 1 289 0 0 0 0 286 38 0 0 2
2727 2344
2743 2344
1 1 288 0 0 0 0 287 39 0 0 2
2696 2344
2712 2344
1 1 287 0 0 0 0 288 40 0 0 2
2661 2344
2677 2344
8 4 291 0 0 4224 0 283 284 0 0 2
2757 2419
2757 2428
7 3 292 0 0 4224 0 283 284 0 0 2
2745 2419
2745 2428
6 2 293 0 0 4224 0 283 284 0 0 2
2733 2419
2733 2428
5 1 294 0 0 4224 0 283 284 0 0 2
2721 2419
2721 2428
0 1 295 0 0 8320 0 0 294 409 0 3
2379 2352
2379 2379
2434 2379
0 2 296 0 0 8320 0 0 294 408 0 4
2418 2352
2418 2367
2446 2367
2446 2379
0 3 297 0 0 12416 0 0 294 407 0 4
2450 2352
2450 2361
2458 2361
2458 2379
4 0 298 0 0 12416 0 294 0 0 406 4
2470 2379
2470 2370
2482 2370
2482 2352
1 1 298 0 0 0 0 292 44 0 0 4
2473 2351
2482 2351
2482 2352
2489 2352
1 1 297 0 0 0 0 291 43 0 0 2
2440 2352
2456 2352
1 1 296 0 0 0 0 290 42 0 0 2
2409 2352
2425 2352
1 1 295 0 0 0 0 289 41 0 0 2
2374 2352
2390 2352
8 4 299 0 0 4224 0 294 293 0 0 2
2470 2427
2470 2436
7 3 300 0 0 4224 0 294 293 0 0 2
2458 2427
2458 2436
6 2 301 0 0 4224 0 294 293 0 0 2
2446 2427
2446 2436
5 1 302 0 0 4224 0 294 293 0 0 2
2434 2427
2434 2436
0 1 303 0 0 8320 0 0 271 421 0 3
2665 2008
2665 2035
2720 2035
0 2 304 0 0 8320 0 0 271 420 0 4
2704 2008
2704 2023
2732 2023
2732 2035
0 3 305 0 0 12416 0 0 271 419 0 4
2736 2008
2736 2017
2744 2017
2744 2035
4 0 306 0 0 12416 0 271 0 0 418 4
2756 2035
2756 2026
2768 2026
2768 2008
1 1 306 0 0 0 0 273 29 0 0 4
2759 2007
2768 2007
2768 2008
2775 2008
1 1 305 0 0 0 0 274 30 0 0 2
2726 2008
2742 2008
1 1 304 0 0 0 0 275 31 0 0 2
2695 2008
2711 2008
1 1 303 0 0 0 0 276 32 0 0 2
2660 2008
2676 2008
8 4 307 0 0 4224 0 271 272 0 0 2
2756 2083
2756 2092
7 3 308 0 0 4224 0 271 272 0 0 2
2744 2083
2744 2092
6 2 309 0 0 4224 0 271 272 0 0 2
2732 2083
2732 2092
5 1 310 0 0 4224 0 271 272 0 0 2
2720 2083
2720 2092
0 1 311 0 0 8320 0 0 282 433 0 3
2378 2016
2378 2043
2433 2043
0 2 312 0 0 8320 0 0 282 432 0 4
2417 2016
2417 2031
2445 2031
2445 2043
0 3 313 0 0 12416 0 0 282 431 0 4
2449 2016
2449 2025
2457 2025
2457 2043
4 0 314 0 0 12416 0 282 0 0 430 4
2469 2043
2469 2034
2481 2034
2481 2016
1 1 314 0 0 0 0 280 36 0 0 4
2472 2015
2481 2015
2481 2016
2488 2016
1 1 313 0 0 0 0 279 35 0 0 2
2439 2016
2455 2016
1 1 312 0 0 0 0 278 34 0 0 2
2408 2016
2424 2016
1 1 311 0 0 0 0 277 33 0 0 2
2373 2016
2389 2016
8 4 315 0 0 4224 0 282 281 0 0 2
2469 2091
2469 2100
7 3 316 0 0 4224 0 282 281 0 0 2
2457 2091
2457 2100
6 2 317 0 0 4224 0 282 281 0 0 2
2445 2091
2445 2100
5 1 318 0 0 4224 0 282 281 0 0 2
2433 2091
2433 2100
0 1 319 0 0 8320 0 0 259 445 0 3
2668 1692
2668 1719
2723 1719
0 2 320 0 0 8320 0 0 259 444 0 4
2707 1692
2707 1707
2735 1707
2735 1719
0 3 321 0 0 12416 0 0 259 443 0 4
2739 1692
2739 1701
2747 1701
2747 1719
4 0 322 0 0 12416 0 259 0 0 442 4
2759 1719
2759 1710
2771 1710
2771 1692
1 1 322 0 0 0 0 261 21 0 0 4
2762 1691
2771 1691
2771 1692
2778 1692
1 1 321 0 0 0 0 262 22 0 0 2
2729 1692
2745 1692
1 1 320 0 0 0 0 263 23 0 0 2
2698 1692
2714 1692
1 1 319 0 0 0 0 264 24 0 0 2
2663 1692
2679 1692
8 4 323 0 0 4224 0 259 260 0 0 2
2759 1767
2759 1776
7 3 324 0 0 4224 0 259 260 0 0 2
2747 1767
2747 1776
6 2 325 0 0 4224 0 259 260 0 0 2
2735 1767
2735 1776
5 1 326 0 0 4224 0 259 260 0 0 2
2723 1767
2723 1776
0 1 327 0 0 8320 0 0 270 457 0 3
2381 1700
2381 1727
2436 1727
0 2 328 0 0 8320 0 0 270 456 0 4
2420 1700
2420 1715
2448 1715
2448 1727
0 3 329 0 0 12416 0 0 270 455 0 4
2452 1700
2452 1709
2460 1709
2460 1727
4 0 330 0 0 12416 0 270 0 0 454 4
2472 1727
2472 1718
2484 1718
2484 1700
1 1 330 0 0 0 0 268 28 0 0 4
2475 1699
2484 1699
2484 1700
2491 1700
1 1 329 0 0 0 0 267 27 0 0 2
2442 1700
2458 1700
1 1 328 0 0 0 0 266 26 0 0 2
2411 1700
2427 1700
1 1 327 0 0 0 0 265 25 0 0 2
2376 1700
2392 1700
8 4 331 0 0 4224 0 270 269 0 0 2
2472 1775
2472 1784
7 3 332 0 0 4224 0 270 269 0 0 2
2460 1775
2460 1784
6 2 333 0 0 4224 0 270 269 0 0 2
2448 1775
2448 1784
5 1 334 0 0 4224 0 270 269 0 0 2
2436 1775
2436 1784
0 1 335 0 0 8320 0 0 306 469 0 3
2658 1070
2658 1097
2713 1097
0 2 336 0 0 8320 0 0 306 468 0 4
2697 1070
2697 1085
2725 1085
2725 1097
0 3 337 0 0 12416 0 0 306 467 0 4
2729 1070
2729 1079
2737 1079
2737 1097
4 0 338 0 0 12416 0 306 0 0 466 4
2749 1097
2749 1088
2761 1088
2761 1070
1 1 338 0 0 0 0 304 52 0 0 4
2752 1069
2761 1069
2761 1070
2768 1070
1 1 337 0 0 0 0 303 51 0 0 2
2719 1070
2735 1070
1 1 336 0 0 0 0 302 50 0 0 2
2688 1070
2704 1070
1 1 335 0 0 0 0 301 49 0 0 2
2653 1070
2669 1070
8 4 339 0 0 4224 0 306 305 0 0 2
2749 1145
2749 1154
7 3 340 0 0 4224 0 306 305 0 0 2
2737 1145
2737 1154
6 2 341 0 0 4224 0 306 305 0 0 2
2725 1145
2725 1154
5 1 342 0 0 4224 0 306 305 0 0 2
2713 1145
2713 1154
0 1 343 0 0 8320 0 0 295 481 0 3
2371 1078
2371 1105
2426 1105
0 2 344 0 0 8320 0 0 295 480 0 4
2410 1078
2410 1093
2438 1093
2438 1105
0 3 345 0 0 12416 0 0 295 479 0 4
2442 1078
2442 1087
2450 1087
2450 1105
4 0 346 0 0 12416 0 295 0 0 478 4
2462 1105
2462 1096
2474 1096
2474 1078
1 1 346 0 0 0 0 297 45 0 0 4
2465 1077
2474 1077
2474 1078
2481 1078
1 1 345 0 0 0 0 298 46 0 0 2
2432 1078
2448 1078
1 1 344 0 0 0 0 299 47 0 0 2
2401 1078
2417 1078
1 1 343 0 0 0 0 300 48 0 0 2
2366 1078
2382 1078
0 1 347 0 0 8320 0 0 318 489 0 3
2657 734
2657 761
2712 761
0 2 348 0 0 8320 0 0 318 488 0 4
2696 734
2696 749
2724 749
2724 761
0 3 349 0 0 12416 0 0 318 487 0 4
2728 734
2728 743
2736 743
2736 761
4 0 350 0 0 12416 0 318 0 0 486 4
2748 761
2748 752
2760 752
2760 734
1 1 350 0 0 0 0 316 60 0 0 4
2751 733
2760 733
2760 734
2767 734
1 1 349 0 0 0 0 315 59 0 0 2
2718 734
2734 734
1 1 348 0 0 0 0 314 58 0 0 2
2687 734
2703 734
1 1 347 0 0 0 0 313 57 0 0 2
2652 734
2668 734
8 4 351 0 0 4224 0 318 317 0 0 2
2748 809
2748 818
7 3 352 0 0 4224 0 318 317 0 0 2
2736 809
2736 818
6 2 353 0 0 4224 0 318 317 0 0 2
2724 809
2724 818
5 1 354 0 0 4224 0 318 317 0 0 2
2712 809
2712 818
0 1 355 0 0 8320 0 0 307 501 0 3
2370 742
2370 769
2425 769
0 2 356 0 0 8320 0 0 307 500 0 4
2409 742
2409 757
2437 757
2437 769
0 3 357 0 0 12416 0 0 307 499 0 4
2441 742
2441 751
2449 751
2449 769
4 0 358 0 0 12416 0 307 0 0 498 4
2461 769
2461 760
2473 760
2473 742
1 1 358 0 0 0 0 309 53 0 0 4
2464 741
2473 741
2473 742
2480 742
1 1 357 0 0 0 0 310 54 0 0 2
2431 742
2447 742
1 1 356 0 0 0 0 311 55 0 0 2
2400 742
2416 742
1 1 355 0 0 0 0 312 56 0 0 2
2365 742
2381 742
8 4 359 0 0 4224 0 307 308 0 0 2
2461 817
2461 826
7 3 360 0 0 4224 0 307 308 0 0 2
2449 817
2449 826
6 2 361 0 0 4224 0 307 308 0 0 2
2437 817
2437 826
5 1 362 0 0 4224 0 307 308 0 0 2
2425 817
2425 826
0 1 363 0 0 8320 0 0 319 513 0 3
2650 151
2650 178
2705 178
0 2 364 0 0 8320 0 0 319 512 0 4
2689 151
2689 166
2717 166
2717 178
0 3 365 0 0 12416 0 0 319 511 0 4
2721 151
2721 160
2729 160
2729 178
4 0 366 0 0 12416 0 319 0 0 510 4
2741 178
2741 169
2753 169
2753 151
1 1 366 0 0 0 0 321 61 0 0 4
2744 150
2753 150
2753 151
2760 151
1 1 365 0 0 0 0 322 62 0 0 2
2711 151
2727 151
1 1 364 0 0 0 0 323 63 0 0 2
2680 151
2696 151
1 1 363 0 0 0 0 324 64 0 0 2
2645 151
2661 151
8 4 367 0 0 4224 0 319 320 0 0 2
2741 226
2741 235
7 3 368 0 0 4224 0 319 320 0 0 2
2729 226
2729 235
6 2 369 0 0 4224 0 319 320 0 0 2
2717 226
2717 235
5 1 370 0 0 4224 0 319 320 0 0 2
2705 226
2705 235
0 1 371 0 0 8320 0 0 331 525 0 3
2363 159
2363 186
2418 186
0 2 372 0 0 8320 0 0 331 524 0 4
2402 159
2402 174
2430 174
2430 186
0 3 373 0 0 12416 0 0 331 523 0 4
2434 159
2434 168
2442 168
2442 186
4 0 374 0 0 12416 0 331 0 0 522 4
2454 186
2454 177
2466 177
2466 159
1 1 374 0 0 0 0 328 68 0 0 4
2457 158
2466 158
2466 159
2473 159
1 1 373 0 0 0 0 327 67 0 0 2
2424 159
2440 159
1 1 372 0 0 0 0 326 66 0 0 2
2393 159
2409 159
1 1 371 0 0 0 0 325 65 0 0 2
2358 159
2374 159
0 1 95 0 0 12416 0 0 350 527 0 4
1294 1736
1269 1736
1269 1820
1374 1820
3 1 95 0 0 0 0 345 349 0 0 3
1271 1695
1294 1695
1294 1771
0 4 375 0 0 8320 0 0 337 529 0 4
1205 1719
1225 1719
1225 2030
1463 2030
3 2 375 0 0 0 0 346 345 0 0 3
1205 1738
1205 1704
1226 1704
8 4 376 0 0 4224 0 331 330 0 0 2
2454 234
2454 243
7 3 377 0 0 4224 0 331 330 0 0 2
2442 234
2442 243
6 2 378 0 0 4224 0 331 330 0 0 2
2430 234
2430 243
5 1 379 0 0 4224 0 331 330 0 0 2
2418 234
2418 243
1 0 380 0 0 4096 0 332 0 0 630 2
486 613
486 614
1 0 3 0 0 0 0 333 0 0 629 2
487 556
487 555
4 0 381 0 0 8320 0 342 0 0 550 3
1589 2061
315 2061
315 522
0 3 380 0 0 4224 0 0 342 551 0 3
305 510
305 2070
1589 2070
2 0 3 0 0 8320 0 342 0 0 552 3
1589 2079
295 2079
295 498
0 1 382 0 0 4224 0 0 342 619 0 3
286 486
286 2088
1589 2088
2 9 383 0 0 8320 0 334 336 0 0 3
214 369
247 369
247 450
1 0 384 0 0 4096 0 335 0 0 542 2
163 368
163 369
1 1 384 0 0 4224 0 334 69 0 0 2
178 369
147 369
0 1 385 0 0 16512 0 0 337 623 0 6
1169 365
1179 365
1179 478
754 478
754 2003
1463 2003
2 0 386 0 0 8320 0 337 0 0 604 6
1463 2012
659 2012
659 832
1188 832
1188 791
1184 791
0 3 387 0 0 16512 0 0 337 583 0 6
1202 1167
1209 1167
1209 1213
664 1213
664 2021
1463 2021
1 0 388 0 0 4096 0 340 0 0 553 2
211 471
211 522
1 0 389 0 0 4096 0 339 0 0 554 2
196 471
196 510
1 0 390 0 0 4096 0 338 0 0 555 2
181 471
181 498
1 0 391 0 0 4096 0 341 0 0 556 2
165 471
165 486
5 0 381 0 0 0 0 336 0 0 618 5
271 522
377 522
377 724
424 724
424 735
0 6 380 0 0 0 0 0 336 630 0 5
427 614
427 596
391 596
391 510
271 510
7 0 3 0 0 0 0 336 0 0 629 3
271 498
423 498
423 555
1 1 388 0 0 8320 0 73 336 0 0 4
148 631
190 631
190 522
223 522
1 2 389 0 0 8320 0 72 336 0 0 4
148 584
180 584
180 510
223 510
1 3 390 0 0 12416 0 71 336 0 0 4
147 538
172 538
172 498
223 498
1 4 391 0 0 4224 0 70 336 0 0 2
147 486
223 486
0 3 381 0 0 0 0 0 350 574 0 3
590 1226
590 1838
1374 1838
3 0 392 0 0 8320 0 349 0 0 575 3
1294 1789
674 1789
674 1154
2 0 393 0 0 4096 0 350 0 0 560 3
1374 1829
692 1829
692 1679
3 2 393 0 0 8320 0 380 349 0 0 4
684 683
692 683
692 1780
1294 1780
0 2 382 0 0 0 0 0 346 576 0 3
737 1126
737 1747
1150 1747
1 4 96 0 0 8320 0 346 343 0 0 4
1150 1729
1145 1729
1145 1603
1132 1603
1 4 97 0 0 4224 0 345 344 0 0 4
1226 1686
989 1686
989 1606
973 1606
4 9 394 0 0 12416 0 349 347 0 0 4
1345 1780
1345 1803
1436 1803
1436 1689
8 4 25 0 0 0 0 348 347 0 0 2
1400 1594
1400 1665
7 3 26 0 0 0 0 348 347 0 0 2
1388 1594
1388 1665
6 2 27 0 0 0 0 348 347 0 0 2
1376 1594
1376 1665
5 1 28 0 0 0 0 348 347 0 0 2
1364 1594
1364 1665
4 9 395 0 0 4224 0 350 352 0 0 3
1425 1829
1626 1829
1626 1689
8 4 9 0 0 0 0 351 352 0 0 2
1590 1597
1590 1665
7 3 10 0 0 0 0 351 352 0 0 2
1578 1597
1578 1665
6 2 11 0 0 0 0 351 352 0 0 2
1566 1597
1566 1665
5 1 12 0 0 0 0 351 352 0 0 2
1554 1597
1554 1665
3 0 381 0 0 0 0 360 0 0 594 5
1369 1296
590 1296
590 1226
578 1226
578 818
0 3 392 0 0 0 0 0 359 595 0 5
653 760
653 1154
674 1154
674 1236
1280 1236
2 0 382 0 0 0 0 356 0 0 599 3
1147 1192
737 1192
737 703
2 0 396 0 0 4224 0 360 0 0 578 3
1369 1287
726 1287
726 1145
3 2 396 0 0 0 0 381 359 0 0 4
684 646
726 646
726 1227
1280 1227
1 0 98 0 0 8320 0 360 0 0 580 3
1369 1278
1262 1278
1262 1140
3 1 98 0 0 0 0 355 359 0 0 3
1259 1140
1280 1140
1280 1218
1 4 100 0 0 8320 0 356 353 0 0 4
1147 1174
1144 1174
1144 1073
1132 1073
1 4 99 0 0 4224 0 355 354 0 0 4
1214 1131
973 1131
973 1070
961 1070
3 2 387 0 0 0 0 356 355 0 0 3
1202 1183
1202 1149
1214 1149
4 9 397 0 0 12416 0 359 357 0 0 4
1331 1227
1331 1266
1429 1266
1429 1157
8 4 29 0 0 0 0 358 357 0 0 2
1393 1074
1393 1133
7 3 30 0 0 0 0 358 357 0 0 2
1381 1074
1381 1133
6 2 31 0 0 0 0 358 357 0 0 2
1369 1074
1369 1133
5 1 32 0 0 0 0 358 357 0 0 2
1357 1074
1357 1133
4 9 398 0 0 8320 0 360 362 0 0 4
1420 1287
1420 1295
1624 1295
1624 1159
8 4 13 0 0 0 0 361 362 0 0 2
1588 1080
1588 1135
7 3 14 0 0 0 0 361 362 0 0 2
1576 1080
1576 1135
6 2 15 0 0 0 0 361 362 0 0 2
1564 1080
1564 1135
5 1 16 0 0 0 0 361 362 0 0 2
1552 1080
1552 1135
3 0 381 0 0 0 0 372 0 0 616 7
1359 887
1340 887
1340 885
578 885
578 818
567 818
567 751
3 0 392 0 0 0 0 367 0 0 617 7
1269 847
1254 847
1254 850
653 850
653 760
638 760
638 735
2 0 399 0 0 4224 0 372 0 0 597 3
1359 878
718 878
718 741
3 2 399 0 0 0 0 382 367 0 0 4
684 600
718 600
718 838
1269 838
2 0 400 0 0 4224 0 384 0 0 624 2
1351 456
689 456
2 0 382 0 0 0 0 363 0 0 619 5
1125 799
737 799
737 703
730 703
730 382
1 0 101 0 0 4224 0 372 0 0 601 3
1359 869
1246 869
1246 758
1 3 101 0 0 0 0 367 364 0 0 4
1269 829
1256 829
1256 758
1237 758
1 4 102 0 0 8320 0 363 366 0 0 4
1125 781
1120 781
1120 696
1108 696
1 4 61 0 0 4224 0 364 365 0 0 4
1192 749
954 749
954 693
939 693
3 2 386 0 0 0 0 363 364 0 0 6
1180 790
1184 790
1184 791
1184 791
1184 767
1192 767
4 9 401 0 0 4224 0 367 369 0 0 4
1320 838
1437 838
1437 750
1420 750
8 4 33 0 0 0 0 368 369 0 0 2
1384 686
1384 726
7 3 34 0 0 0 0 368 369 0 0 2
1372 686
1372 726
6 2 35 0 0 0 0 368 369 0 0 2
1360 686
1360 726
5 1 36 0 0 0 0 368 369 0 0 2
1348 686
1348 726
4 9 402 0 0 4224 0 372 370 0 0 3
1410 878
1619 878
1619 751
8 4 17 0 0 0 0 371 370 0 0 2
1583 685
1583 727
7 3 18 0 0 0 0 371 370 0 0 2
1571 685
1571 727
6 2 19 0 0 0 0 371 370 0 0 2
1559 685
1559 727
5 1 20 0 0 0 0 371 370 0 0 2
1547 685
1547 727
0 1 103 0 0 8320 0 0 384 621 0 3
1245 356
1245 447
1351 447
3 0 381 0 0 0 0 384 0 0 618 5
1351 465
713 465
713 751
560 751
560 735
2 3 392 0 0 0 0 377 385 0 0 6
633 735
708 735
708 418
1256 418
1256 417
1265 417
0 1 381 0 0 0 0 0 377 0 0 2
415 735
597 735
8 2 382 0 0 0 0 336 376 0 0 6
271 486
412 486
412 490
526 490
526 382
1114 382
1 4 104 0 0 8320 0 376 373 0 0 4
1114 364
1112 364
1112 302
1099 302
1 3 103 0 0 0 0 385 375 0 0 4
1265 399
1258 399
1258 356
1233 356
1 4 62 0 0 4224 0 375 374 0 0 4
1188 347
947 347
947 295
926 295
3 2 385 0 0 0 0 376 375 0 0 3
1169 373
1169 365
1188 365
2 3 400 0 0 0 0 385 383 0 0 4
1265 408
689 408
689 564
684 564
0 1 3 0 0 0 0 0 380 629 0 3
533 555
533 674
639 674
0 2 380 0 0 0 0 0 380 627 0 3
523 626
523 692
639 692
2 0 380 0 0 0 0 382 0 0 630 5
639 609
611 609
611 626
523 626
523 614
1 0 403 0 0 8192 0 382 0 0 632 3
639 591
619 591
619 555
0 1 3 0 0 0 0 0 379 0 0 2
413 555
550 555
0 1 380 0 0 0 0 0 378 0 0 2
414 614
549 614
2 2 2 0 0 0 0 383 378 0 0 3
639 573
585 573
585 614
1 2 403 0 0 4224 0 383 379 0 0 2
639 555
586 555
4 9 404 0 0 4224 0 384 389 0 0 3
1402 456
1613 456
1613 338
4 9 405 0 0 8320 0 385 387 0 0 5
1316 408
1316 417
1430 417
1430 331
1416 331
8 4 21 0 0 0 0 388 389 0 0 2
1577 280
1577 314
7 3 22 0 0 0 0 388 389 0 0 2
1565 280
1565 314
6 2 23 0 0 0 0 388 389 0 0 2
1553 280
1553 314
5 1 24 0 0 0 0 388 389 0 0 2
1541 280
1541 314
8 4 37 0 0 0 0 386 387 0 0 2
1380 275
1380 307
7 3 38 0 0 0 0 386 387 0 0 2
1368 275
1368 307
6 2 39 0 0 0 0 386 387 0 0 2
1356 275
1356 307
5 1 40 0 0 0 0 386 387 0 0 2
1344 275
1344 307
19
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 6
26 511 94 534
38 521 81 536
6 LINHAS
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 4
29 615 84 638
42 625 70 640
4 BYTE
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
38 466 84 489
50 476 71 491
3 TAG
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 8
1518 37 1603 61
1528 45 1592 61
8 BYTE = 1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 8
1323 34 1408 58
1333 42 1397 58
8 BYTE = 0
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
1039 216 1084 240
1049 224 1073 240
3 TAG
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
879 215 924 239
889 223 913 239
3 USO
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 196
39 18 284 262
49 26 273 218
196 Cache 4 linhas com 2 colunas 
cada de uma de 4 bits

Memoria principal
16 linhas de 4 bits
8 conj's pois s�o 2 colunas 
na cache

MAPEAMENTO DIRETO

USO TAG LINHA BYTE
 1   1    2    1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
2396 75 2441 99
2406 83 2430 99
3 PAR
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 5
2674 69 2735 93
2684 77 2724 93
5 IMPAR
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 10
2535 2416 2636 2440
2545 2424 2625 2440
10 CONJUNTO 7
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 10
2518 198 2619 222
2528 206 2608 222
10 CONJUNTO 0
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 10
2518 488 2619 512
2528 496 2608 512
10 CONJUNTO 1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 10
2516 774 2617 798
2526 782 2606 798
10 CONJUNTO 2
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 10
2521 1142 2622 1166
2531 1150 2611 1166
10 CONJUNTO 3
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 10
2521 1440 2622 1464
2531 1448 2611 1464
10 CONJUNTO 4
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 10
2537 1746 2638 1770
2547 1754 2627 1770
10 CONJUNTO 5
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 10
2538 2072 2639 2096
2548 2080 2628 2096
10 CONJUNTO 6
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 146
240 143 581 247
250 151 570 231
146 A tag s� ser� recebida se der miss e ele 
selecinar o conjunto x, a partir de x 
ele define se � tag 0 ou 1:
conjunto 0-3: 0
conjunto 4-7: 1
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0

CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 1050 1 90 10
176 80 1918 1019
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
2 4 0.500000 0.500000
344 176 457 273
42991634 0
0
6 Title:
5 Name:
0
0
0
554
13 Logic Switch~
5 134 1051 0 1 11
0 9
0
0 0 21344 0
2 0V
-32 -4 -18 4
4 Auto
-40 -13 -12 -5
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
5130 0 0
2
44286.3 0
0
13 Logic Switch~
5 2699 482 0 10 11
0 83 0 0 0 0 0 0 0 0
1
0
0 0 21344 0
2 5V
-32 -4 -18 4
3 V14
-34 -17 -13 -9
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
391 0 0
2
5.89979e-315 0
0
13 Logic Switch~
5 2400 487 0 10 11
0 84 0 0 0 0 0 0 0 0
1
0
0 0 21344 0
2 5V
-32 -4 -18 4
3 V13
-34 -17 -13 -9
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
3124 0 0
2
5.89979e-315 5.26354e-315
0
13 Logic Switch~
5 2084 499 0 10 11
0 85 0 0 0 0 0 0 0 0
1
0
0 0 21344 0
2 5V
-32 -4 -18 4
2 V6
-31 -17 -17 -9
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
3421 0 0
2
5.89979e-315 5.30499e-315
0
13 Logic Switch~
5 1862 499 0 10 11
0 87 0 0 0 0 0 0 0 0
1
0
0 0 21344 0
2 5V
-32 -4 -18 4
3 V15
-34 -17 -13 -9
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
8157 0 0
2
5.89979e-315 5.32571e-315
0
13 Logic Switch~
5 1722 558 0 1 11
0 89
0
0 0 21344 0
2 0V
-32 -4 -18 4
7 Vlibera
-48 -17 1 -9
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
5572 0 0
2
5.89979e-315 5.34643e-315
0
13 Logic Switch~
5 599 1162 0 10 11
0 92 0 0 0 0 0 0 0 0
1
0
0 0 21344 0
2 5V
-32 -4 -18 4
6 Manual
-47 -13 -5 -5
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
8901 0 0
2
5.89979e-315 5.3568e-315
0
13 Logic Switch~
5 219 893 0 1 11
0 40
0
0 0 21344 0
2 0V
-6 -16 8 -8
5 Reset
-16 -26 19 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
7361 0 0
2
44286.3 1
0
13 Logic Switch~
5 782 1613 0 1 11
0 346
0
0 0 21344 0
2 0V
-6 -16 8 -8
5 Vbit1
-17 -26 18 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
4747 0 0
2
5.89979e-315 5.36716e-315
0
13 Logic Switch~
5 780 1557 0 1 11
0 345
0
0 0 21344 0
2 0V
-6 -16 8 -8
5 Vbit2
-17 -26 18 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
972 0 0
2
5.89979e-315 5.37752e-315
0
13 Logic Switch~
5 1159 1677 0 1 11
0 343
0
0 0 21344 0
2 0V
-6 -16 8 -8
3 V32
-10 -26 11 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3472 0 0
2
44286.3 2
0
13 Logic Switch~
5 1260 1570 0 10 11
0 412 0 0 0 0 0 0 0 0
1
0
0 0 21344 270
2 5V
-6 -21 8 -13
3 V29
-10 -31 11 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
9998 0 0
2
5.89979e-315 5.38788e-315
0
13 Logic Switch~
5 1357 1567 0 10 11
0 411 0 0 0 0 0 0 0 0
1
0
0 0 21344 270
2 5V
-6 -21 8 -13
3 V22
-10 -31 11 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
3536 0 0
2
5.89979e-315 5.39306e-315
0
13 Logic Switch~
5 1440 1566 0 10 11
0 410 0 0 0 0 0 0 0 0
1
0
0 0 21344 270
2 5V
-6 -21 8 -13
3 V30
-10 -31 11 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
4597 0 0
2
5.89979e-315 5.39824e-315
0
13 Logic Switch~
5 1528 1573 0 10 11
0 409 0 0 0 0 0 0 0 0
1
0
0 0 21344 270
2 5V
-6 -21 8 -13
3 V31
-10 -31 11 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
3835 0 0
2
5.89979e-315 5.40342e-315
0
13 Logic Switch~
5 822 970 0 1 11
0 414
0
0 0 21344 270
2 0V
-6 -21 8 -13
3 V28
-9 -31 12 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3670 0 0
2
5.89979e-315 5.4086e-315
0
13 Logic Switch~
5 859 970 0 1 11
0 413
0
0 0 21344 270
2 0V
-6 -21 8 -13
3 V11
-9 -31 12 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
5616 0 0
2
5.89979e-315 5.41378e-315
0
13 Logic Switch~
5 783 970 0 1 11
0 415
0
0 0 21344 270
2 0V
-6 -21 8 -13
3 V10
-9 -31 12 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
9323 0 0
2
5.89979e-315 5.41896e-315
0
13 Logic Switch~
5 746 970 0 1 11
0 416
0
0 0 21344 270
2 0V
-6 -21 8 -13
2 V8
-6 -31 8 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
317 0 0
2
5.89979e-315 5.42414e-315
0
13 Logic Switch~
5 317 1748 0 10 11
0 421 0 0 0 0 0 0 0 0
1
0
0 0 21344 0
2 5V
-6 -16 8 -8
4 SET1
-12 -26 16 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
3108 0 0
2
5.89979e-315 5.42933e-315
0
13 Logic Switch~
5 1306 1025 0 1 11
0 156
0
0 0 21344 270
2 0V
-6 -21 8 -13
2 VE
-7 -31 7 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
4299 0 0
2
44286.3 3
0
13 Logic Switch~
5 1285 1025 0 10 11
0 155 0 0 0 0 0 0 0 0
1
0
0 0 21344 270
2 5V
-6 -21 8 -13
3 VEL
-10 -31 11 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
9672 0 0
2
44286.3 4
0
8 2-In OR~
219 876 1395 0 3 22
0 4 3 2
0
0 0 608 0
6 74LS32
-21 -24 21 -16
5 U182B
-10 -25 25 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 91 0
1 U
7876 0 0
2
44286.3 5
0
8 3-In OR~
219 1276 798 0 4 22
0 5 6 7 27
0
0 0 608 270
4 4075
-14 -24 14 -16
5 U177C
0 -4 35 4
0
15 DVDD=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 11 12 13 10 3 4 5 6 1
2 8 9 11 12 13 10 0 0 0
0 1 0
65 0 0 0 3 3 82 0
1 U
6369 0 0
2
44286.3 6
0
10 Buffer 3S~
219 774 614 0 3 22
0 10 9 11
0
0 0 608 0
8 BUFFER3S
-27 -51 29 -43
5 U178D
-18 -20 17 -12
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
0
22

0 12 13 11 2 1 3 5 4 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 84 0
1 U
9172 0 0
2
44286.3 7
0
9 Inverter~
13 707 616 0 2 22
0 12 10
0
0 0 608 692
6 74LS04
-21 -19 21 -11
5 U184C
-18 -20 17 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 5 6 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 3 89 0
1 U
7100 0 0
2
44286.3 8
0
5 4082~
219 1354 738 0 5 22
0 22 21 19 20 8
0
0 0 608 270
4 4082
-7 -24 21 -16
5 U174B
-17 -12 18 -4
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
13 type: digital
5 DIP14
22

0 9 10 11 12 13 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 0 2 2 90 0
1 U
3820 0 0
2
44286.3 9
0
8 2-In OR~
219 1170 782 0 3 22
0 28 29 30
0
0 0 608 270
6 74LS32
-21 -24 21 -16
5 U182A
-14 -3 21 5
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 91 0
1 U
7678 0 0
2
44286.3 10
0
8 2-In OR~
219 1101 782 0 3 22
0 32 33 31
0
0 0 608 270
6 74LS32
-21 -24 21 -16
5 U179D
-14 -3 21 5
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 85 0
1 U
961 0 0
2
44286.3 11
0
5 4082~
219 1281 738 0 5 22
0 22 21 23 20 6
0
0 0 608 270
4 4082
-7 -24 21 -16
5 U173B
-17 -12 18 -4
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
13 type: digital
5 DIP14
22

0 9 10 11 12 13 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 0 2 2 88 0
1 U
3178 0 0
2
44286.3 12
0
5 4082~
219 1243 738 0 5 22
0 22 21 23 24 7
0
0 0 608 270
4 4082
-7 -24 21 -16
5 U174A
-17 -12 18 -4
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
13 type: digital
5 DIP14
22

0 2 3 4 5 1 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 0 2 1 90 0
1 U
3409 0 0
2
44286.3 13
0
5 4082~
219 1205 738 0 5 22
0 26 25 19 20 28
0
0 0 608 270
4 4082
-7 -24 21 -16
5 U173A
-17 -12 18 -4
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
13 type: digital
5 DIP14
22

0 2 3 4 5 1 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 0 2 1 88 0
1 U
3951 0 0
2
44286.3 14
0
5 4082~
219 1130 738 0 5 22
0 26 25 23 20 32
0
0 0 608 270
4 4082
-7 -24 21 -16
5 U154B
-17 -12 18 -4
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
13 type: digital
5 DIP14
22

0 9 10 11 12 13 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 0 2 2 79 0
1 U
8885 0 0
2
44286.3 15
0
5 4082~
219 1094 738 0 5 22
0 26 25 23 24 33
0
0 0 608 270
4 4082
-7 -24 21 -16
4 U63A
-14 -12 14 -4
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
13 type: digital
5 DIP14
22

0 2 3 4 5 1 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 0 2 1 78 0
1 U
3780 0 0
2
44286.3 16
0
5 4082~
219 1318 738 0 5 22
0 22 21 19 24 5
0
0 0 608 270
4 4082
-7 -24 21 -16
5 U154A
-17 -12 18 -4
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
13 type: digital
5 DIP14
22

0 2 3 4 5 1 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 0 2 1 79 0
1 U
9265 0 0
2
44286.3 17
0
5 4082~
219 1168 738 0 5 22
0 26 25 19 24 29
0
0 0 608 270
4 4082
-7 -24 21 -16
4 U63B
-14 -12 14 -4
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
13 type: digital
5 DIP14
22

0 9 10 11 12 13 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 0 2 2 78 0
1 U
9442 0 0
2
44286.3 18
0
5 4082~
219 1059 738 0 5 22
0 26 21 19 20 35
0
0 0 608 270
4 4082
-7 -24 21 -16
4 U37A
-14 -12 14 -4
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
13 type: digital
5 DIP14
22

0 2 3 4 5 1 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 0 2 1 65 0
1 U
9424 0 0
2
44286.3 19
0
9 Inverter~
13 939 614 0 2 22
0 22 26
0
0 0 608 0
6 74LS04
-21 -19 21 -11
5 U184B
-14 -13 21 -5
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 3 4 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 2 89 0
1 U
9968 0 0
2
44286.3 20
0
5 4082~
219 1025 738 0 5 22
0 26 21 19 24 34
0
0 0 608 270
4 4082
-7 -24 21 -16
4 U28B
-14 -12 14 -4
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
13 type: digital
5 DIP14
22

0 9 10 11 12 13 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 0 2 2 7 0
1 U
9281 0 0
2
44286.3 21
0
5 4082~
219 990 738 0 5 22
0 26 21 23 20 36
0
0 0 608 270
4 4082
-7 -24 21 -16
4 U28A
-14 -12 14 -4
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
13 type: digital
5 DIP14
22

0 2 3 4 5 1 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 0 2 1 7 0
1 U
8464 0 0
2
44286.3 22
0
5 4082~
219 955 738 0 5 22
0 26 21 23 24 37
0
0 0 608 270
4 4082
-7 -24 21 -16
3 U8B
-11 -12 10 -4
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
13 type: digital
5 DIP14
22

0 9 10 11 12 13 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 0 2 2 3 0
1 U
7168 0 0
2
44286.3 23
0
8 4-In OR~
219 983 798 0 5 22
0 35 34 36 37 38
0
0 0 608 270
4 4072
-14 -24 14 -16
3 U9A
-9 -5 12 3
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
12 type:digital
5 DIP14
22

0 2 3 4 5 1 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 0 2 1 4 0
1 U
3171 0 0
2
44286.3 24
0
8 2-In OR~
219 642 613 0 3 22
0 40 8 12
0
0 0 608 692
6 74LS32
-21 -24 21 -16
5 U179C
-10 -25 25 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 9 10 8 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 85 0
1 U
4139 0 0
2
44286.3 25
0
10 Buffer 3S~
219 889 212 0 3 22
0 43 9 22
0
0 0 608 0
8 BUFFER3S
-27 -51 29 -43
5 U178C
-18 -20 17 -12
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
0
22

0 9 10 8 2 1 3 5 4 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 84 0
1 U
6435 0 0
2
44286.3 26
0
14 Logic Display~
6 809 183 0 1 2
10 43
0
0 0 53872 512
6 100MEG
3 -16 45 -8
4 L163
-14 -21 14 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
5283 0 0
2
44286.3 27
0
12 D Flip-Flop~
219 778 248 0 4 9
0 41 18 612 43
0
0 0 4704 0
3 DFF
-10 -53 11 -45
2 U5
-7 -55 7 -47
0
14 DVCC=6;DGND=5;
47 %D [%6bi %5bi %1i %2i][%6bo %1o %2o %3o %4o] %M
0
11 typeDigital
4 DIP6
9

0 1 2 3 4 1 2 3 4 0
65 0 0 512 1 0 0 0
1 U
6874 0 0
2
44286.3 28
0
8 4-In OR~
219 945 892 0 5 22
0 50 38 92 613 39
0
0 0 608 0
4 4072
-14 -24 14 -16
3 U4A
2 -11 23 -3
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
12 type:digital
5 DIP14
22

0 2 3 4 5 1 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 512 2 1 2 0
1 U
5305 0 0
2
5.89979e-315 5.43192e-315
0
13 Quad 3-State~
48 1010 536 0 9 19
0 44 45 46 43 49 48 47 42 12
0
0 0 4704 0
8 QUAD3STA
-28 -44 28 -36
2 U3
-7 -46 7 -38
0
15 DVCC=16;DGND=8;
85 %D [%16bi %8bi %1i %2i %3i %4i %9i]
+ [%16bo %1o %2o %3o %4o %9o %5o %6o %7o %8o] %M
0
12 type:digital
5 DIP16
19

0 1 2 3 4 5 6 7 8 9
1 2 3 4 5 6 7 8 9 0
65 0 0 0 1 0 0 0
1 U
34 0 0
2
44286.3 29
0
5 4073~
219 260 1619 0 4 22
0 71 51 3 54
0
0 0 608 512
4 4073
-7 -24 21 -16
5 U175B
-20 -25 15 -17
0
15 DVDD=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 1 2 8 9 3 4 5 6 1
2 8 9 11 12 13 10 0 0 0
0 1 0
65 0 0 0 3 2 80 0
1 U
969 0 0
2
44286.3 30
0
9 Inverter~
13 358 1787 0 2 22
0 53 52
0
0 0 608 0
6 74LS04
-21 -19 21 -11
3 z2D
-7 -9 14 -1
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 9 8 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 4 73 0
1 U
8402 0 0
2
44286.3 31
0
5 4071~
219 311 1807 0 3 22
0 9 614 53
0
0 0 608 0
4 4071
-7 -24 21 -16
5 U185A
-11 -15 24 -7
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 512 4 1 86 0
1 U
3751 0 0
2
44286.3 32
0
13 Quad 3-State~
48 346 1055 0 9 19
0 58 57 56 55 66 65 64 63 54
0
0 0 4704 0
8 QUAD3STA
-28 -44 28 -36
4 U180
-14 -46 14 -38
0
15 DVCC=16;DGND=8;
85 %D [%16bi %8bi %1i %2i %3i %4i %9i]
+ [%16bo %1o %2o %3o %4o %9o %5o %6o %7o %8o] %M
0
12 type:digital
5 DIP16
19

0 1 2 3 4 5 6 7 8 9
1 2 3 4 5 6 7 8 9 0
65 0 0 0 1 0 0 0
1 U
4292 0 0
2
44286.3 33
0
9 Inverter~
13 211 1604 0 2 22
0 54 72
0
0 0 608 602
6 74LS04
-21 -19 21 -11
5 U184A
-18 0 17 8
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 1 89 0
1 U
6118 0 0
2
44286.3 34
0
13 Quad 3-State~
48 214 1540 0 9 19
0 67 68 69 70 62 61 60 59 72
0
0 0 4704 512
8 QUAD3STA
-28 -44 28 -36
4 U183
-14 -46 14 -38
0
15 DVCC=16;DGND=8;
85 %D [%16bi %8bi %1i %2i %3i %4i %9i]
+ [%16bo %1o %2o %3o %4o %9o %5o %6o %7o %8o] %M
0
12 type:digital
5 DIP16
19

0 1 2 3 4 5 6 7 8 9
1 2 3 4 5 6 7 8 9 0
65 0 0 0 1 0 0 0
1 U
34 0 0
2
44286.3 35
0
5 4071~
219 453 1136 0 3 22
0 63 59 73
0
0 0 608 0
4 4071
-7 -24 21 -16
5 U181D
-5 -11 30 -3
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 4 87 0
1 U
6357 0 0
2
44286.3 36
0
5 4071~
219 453 1102 0 3 22
0 64 60 74
0
0 0 608 0
4 4071
-7 -24 21 -16
5 U181C
-5 -11 30 -3
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 8 9 10 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 3 87 0
1 U
319 0 0
2
44286.3 37
0
5 4071~
219 454 1068 0 3 22
0 65 61 75
0
0 0 608 0
4 4071
-7 -24 21 -16
5 U181B
-5 -11 30 -3
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 5 6 4 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 2 87 0
1 U
3976 0 0
2
44286.3 38
0
5 4071~
219 455 1034 0 3 22
0 66 62 76
0
0 0 608 0
4 4071
-7 -24 21 -16
5 U181A
-5 -11 30 -3
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 1 87 0
1 U
7634 0 0
2
44286.3 39
0
5 4025~
219 657 1405 0 4 22
0 71 78 102 50
0
0 0 608 0
4 4025
-14 -24 14 -16
5 U143A
-10 -25 25 -17
0
15 DVDD=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 3 4 5 6 3 4 5 6 1
2 8 9 11 12 13 10 0 0 0
0 2 0
65 0 0 0 3 1 57 0
1 U
523 0 0
2
44286.3 40
0
9 2-In AND~
219 1635 1536 0 3 22
0 78 3 17
0
0 0 608 0
6 74LS08
-21 -24 21 -16
5 U166D
-19 -25 16 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 69 0
1 U
6748 0 0
2
5.89979e-315 5.43451e-315
0
10 Buffer 3S~
219 2731 482 0 3 22
0 83 79 80
0
0 0 608 0
8 BUFFER3S
-27 -51 29 -43
5 U178B
-18 -20 17 -12
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
0
22

0 5 4 6 2 1 3 5 4 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 84 0
1 U
6901 0 0
2
5.89979e-315 5.4371e-315
0
10 Buffer 3S~
219 2432 487 0 3 22
0 84 79 81
0
0 0 608 0
8 BUFFER3S
-27 -51 29 -43
5 U178A
-18 -20 17 -12
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
0
22

0 2 1 3 2 1 3 5 4 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 84 0
1 U
842 0 0
2
5.89979e-315 5.43969e-315
0
10 Buffer 3S~
219 2116 499 0 3 22
0 85 79 82
0
0 0 608 0
8 BUFFER3S
-27 -51 29 -43
5 U167D
-18 -20 17 -12
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
0
22

0 12 13 11 2 1 3 5 4 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 83 0
1 U
3277 0 0
2
5.89979e-315 5.44228e-315
0
10 Buffer 3S~
219 1894 499 0 3 22
0 87 79 86
0
0 0 608 0
8 BUFFER3S
-27 -51 29 -43
5 U167C
-18 -20 17 -12
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
0
22

0 9 10 8 2 1 3 5 4 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 83 0
1 U
4212 0 0
2
5.89979e-315 5.44487e-315
0
9 Inverter~
13 1693 635 0 2 22
0 17 79
0
0 0 608 692
6 74LS04
-21 -19 21 -11
3 z5F
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 13 12 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 6 77 0
1 U
4720 0 0
2
5.89979e-315 5.44746e-315
0
10 Buffer 3S~
219 1754 558 0 3 22
0 89 79 88
0
0 0 608 0
8 BUFFER3S
-27 -51 29 -43
5 U167B
-18 -20 17 -12
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
0
22

0 5 4 6 2 1 3 5 4 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 83 0
1 U
5551 0 0
2
5.89979e-315 5.45005e-315
0
8 2-In OR~
219 2770 542 0 3 22
0 16 80 91
0
0 0 608 270
6 74LS32
-21 -24 21 -16
5 U141A
-11 -3 24 5
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 56 0
1 U
6986 0 0
2
5.89979e-315 5.45264e-315
0
8 2-In OR~
219 2469 537 0 3 22
0 15 81 606
0
0 0 608 270
6 74LS32
-21 -24 21 -16
5 U171D
-11 -3 24 5
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 76 0
1 U
8745 0 0
2
5.89979e-315 5.45523e-315
0
8 2-In OR~
219 2171 536 0 3 22
0 14 82 605
0
0 0 608 270
6 74LS32
-21 -24 21 -16
5 U171C
-11 -6 24 2
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 9 10 8 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 76 0
1 U
9592 0 0
2
5.89979e-315 5.45782e-315
0
8 2-In OR~
219 1812 598 0 3 22
0 17 88 90
0
0 0 608 270
6 74LS32
-21 -24 21 -16
5 U171B
-11 -3 24 5
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 76 0
1 U
8748 0 0
2
5.89979e-315 5.46041e-315
0
8 2-In OR~
219 1959 530 0 3 22
0 13 86 607
0
0 0 608 270
6 74LS32
-21 -24 21 -16
5 U171B
-11 -3 24 5
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 76 0
1 U
7168 0 0
2
5.89979e-315 5.463e-315
0
8 3-In OR~
219 1041 1986 0 4 22
0 197 193 218 400
0
0 0 608 270
4 4075
-14 -24 14 -16
5 U177B
-10 -6 25 2
0
15 DVDD=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 1 2 8 9 3 4 5 6 1
2 8 9 11 12 13 10 0 0 0
0 1 0
65 0 0 0 3 2 82 0
1 U
631 0 0
2
44286.3 41
0
8 3-In OR~
219 1004 1988 0 4 22
0 196 192 219 399
0
0 0 608 270
4 4075
-14 -24 14 -16
5 U177A
-10 -6 25 2
0
15 DVDD=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 3 4 5 6 3 4 5 6 1
2 8 9 11 12 13 10 0 0 0
0 1 0
65 0 0 0 3 1 82 0
1 U
9466 0 0
2
44286.3 42
0
8 3-In OR~
219 968 1989 0 4 22
0 195 191 220 398
0
0 0 608 270
4 4075
-14 -24 14 -16
5 U176C
-10 -6 25 2
0
15 DVDD=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 11 12 13 10 3 4 5 6 1
2 8 9 11 12 13 10 0 0 0
0 1 0
65 0 0 0 3 3 81 0
1 U
3266 0 0
2
44286.3 43
0
8 3-In OR~
219 928 1987 0 4 22
0 194 190 221 397
0
0 0 608 270
4 4075
-14 -24 14 -16
5 U176B
-10 -6 25 2
0
15 DVDD=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 1 2 8 9 3 4 5 6 1
2 8 9 11 12 13 10 0 0 0
0 1 0
65 0 0 0 3 2 81 0
1 U
7693 0 0
2
44286.3 44
0
13 Quad 3-State~
48 1128 965 0 9 19
0 100 99 98 97 96 95 94 93 101
0
0 0 4704 692
8 QUAD3STA
-28 -44 28 -36
4 U164
-14 46 14 54
0
15 DVCC=16;DGND=8;
85 %D [%16bi %8bi %1i %2i %3i %4i %9i]
+ [%16bo %1o %2o %3o %4o %9o %5o %6o %7o %8o] %M
0
12 type:digital
5 DIP16
19

0 1 2 3 4 5 6 7 8 9
1 2 3 4 5 6 7 8 9 0
65 0 0 0 1 0 0 0
1 U
3723 0 0
2
44286.3 45
0
9 Inverter~
13 1125 916 0 2 22
0 39 101
0
0 0 608 270
6 74LS04
-21 -19 21 -11
3 z5E
16 -8 37 0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 11 10 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 5 77 0
1 U
3440 0 0
2
44286.3 46
0
9 Inverter~
13 890 1358 0 2 22
0 31 103
0
0 0 608 0
6 74LS04
-21 -19 21 -11
3 z5D
-10 -3 11 5
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 9 8 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 4 77 0
1 U
6263 0 0
2
44286.3 47
0
10 Buffer 3S~
219 1310 1409 0 3 22
0 132 30 133
0
0 0 608 692
8 BUFFER3S
-27 -51 29 -43
5 U167A
-18 14 17 22
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
0
22

0 2 1 3 2 1 3 5 4 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 83 0
1 U
4900 0 0
2
44286.3 48
0
13 Quad 3-State~
48 1224 1345 0 9 19
0 104 105 106 107 111 110 109 108 103
0
0 0 4704 0
8 QUAD3STA
-28 -44 28 -36
4 U157
-14 -46 14 -38
0
15 DVCC=16;DGND=8;
85 %D [%16bi %8bi %1i %2i %3i %4i %9i]
+ [%16bo %1o %2o %3o %4o %9o %5o %6o %7o %8o] %M
0
12 type:digital
5 DIP16
19

0 1 2 3 4 5 6 7 8 9
1 2 3 4 5 6 7 8 9 0
65 0 0 0 1 0 0 0
1 U
8783 0 0
2
44286.3 49
0
10 Buffer 3S~
219 959 1168 0 3 22
0 132 39 112
0
0 0 608 90
8 BUFFER3S
-27 -51 29 -43
5 U139A
-49 -5 -14 3
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
0
22

0 2 1 3 2 1 3 5 4 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 58 0
1 U
3221 0 0
2
44286.3 50
0
12 Quad D Flop~
47 959 1086 0 9 19
0 126 125 124 123 100 99 98 97 112
0
0 0 4704 0
4 QDFF
-14 -44 14 -36
2 U1
-8 -46 6 -38
0
15 DVCC=16;DGND=8;
85 %D [%16bi %8bi %1i %2i %3i %4i %9i]
+ [%16bo %1o %2o %3o %4o %9o %5o %6o %7o %8o] %M
0
11 typeDigital
5 DIP16
19

0 1 2 3 4 5 6 7 8 9
1 2 3 4 5 6 7 8 9 0
65 0 0 0 1 0 0 0
1 U
3215 0 0
2
44286.3 51
0
10 Buffer 3S~
219 574 814 0 3 22
0 8 9 113
0
0 0 608 512
8 BUFFER3S
-27 -51 29 -43
5 U168B
-18 -20 17 -12
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
0
22

0 5 4 6 2 1 3 5 4 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 71 0
1 U
7903 0 0
2
44286.3 52
0
10 Buffer 3S~
219 414 837 0 3 22
0 50 113 115
0
0 0 608 90
8 BUFFER3S
-27 -51 29 -43
1 k
-3 -3 4 5
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
0
22

0 2 1 3 2 1 3 5 4 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 72 0
1 U
7121 0 0
2
44286.3 53
0
10 Buffer 3S~
219 381 836 0 3 22
0 114 113 116
0
0 0 608 90
8 BUFFER3S
-27 -51 29 -43
1 g
-4 -1 3 7
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
0
22

0 2 1 3 2 1 3 5 4 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 70 0
1 U
4484 0 0
2
44286.3 54
0
9 2-In AND~
219 788 1342 0 3 22
0 31 51 117
0
0 0 608 0
6 74LS08
-21 -24 21 -16
5 U166C
-11 -13 24 -5
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 69 0
1 U
5996 0 0
2
44286.3 55
0
9 Inverter~
13 934 643 0 2 22
0 25 21
0
0 0 608 0
6 74LS04
-21 -19 21 -11
3 z5C
-11 -6 10 2
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 5 6 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 3 77 0
1 U
7804 0 0
2
44286.3 56
0
9 Inverter~
13 926 669 0 2 22
0 19 23
0
0 0 608 0
6 74LS04
-21 -19 21 -11
3 z5B
-11 -6 10 2
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 3 4 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 2 77 0
1 U
5523 0 0
2
44286.3 57
0
14 Logic Display~
6 813 288 0 1 2
10 46
0
0 0 53872 512
6 100MEG
3 -16 45 -8
4 L162
-14 -21 14 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3330 0 0
2
44286.3 58
0
10 Buffer 3S~
219 890 321 0 3 22
0 46 9 25
0
0 0 608 0
8 BUFFER3S
-27 -51 29 -43
5 U170D
-18 -20 17 -12
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
0
22

0 12 13 11 2 1 3 5 4 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 75 0
1 U
3465 0 0
2
44286.3 59
0
12 D Flip-Flop~
219 780 357 0 4 9
0 118 18 615 46
0
0 0 4704 0
3 DFF
-10 -53 11 -45
4 U172
-14 -55 14 -47
0
14 DVCC=6;DGND=5;
47 %D [%6bi %5bi %1i %2i][%6bo %1o %2o %3o %4o] %M
0
11 typeDigital
4 DIP6
9

0 1 2 3 4 1 2 3 4 0
65 0 0 512 1 0 0 0
1 U
8396 0 0
2
44286.3 60
0
9 2-In AND~
219 788 1422 0 3 22
0 27 51 3
0
0 0 608 0
6 74LS08
-21 -24 21 -16
5 U166B
-11 -13 24 -5
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 69 0
1 U
3685 0 0
2
44286.3 61
0
9 2-In AND~
219 788 1380 0 3 22
0 30 51 4
0
0 0 608 0
6 74LS08
-21 -24 21 -16
5 U166A
-11 -13 24 -5
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 69 0
1 U
7849 0 0
2
5.89979e-315 5.46559e-315
0
14 Logic Display~
6 1268 910 0 1 2
10 122
0
0 0 53872 512
6 100MEG
3 -16 45 -8
3 L50
-11 -21 10 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
6343 0 0
2
5.89979e-315 5.46818e-315
0
14 Logic Display~
6 1245 910 0 1 2
10 121
0
0 0 53872 512
6 100MEG
3 -16 45 -8
3 L51
-11 -21 10 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
7376 0 0
2
5.89979e-315 5.47077e-315
0
14 Logic Display~
6 1223 910 0 1 2
10 120
0
0 0 53872 512
6 100MEG
3 -16 45 -8
3 L52
-11 -21 10 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
9156 0 0
2
5.89979e-315 5.47207e-315
0
14 Logic Display~
6 1201 910 0 1 2
10 119
0
0 0 53872 512
6 100MEG
3 -16 45 -8
3 L55
-11 -21 10 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
5776 0 0
2
5.89979e-315 5.47336e-315
0
14 Logic Display~
6 940 937 0 1 2
10 126
0
0 0 53872 512
6 100MEG
3 -16 45 -8
4 L161
-14 -21 14 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
7207 0 0
2
5.89979e-315 5.47466e-315
0
14 Logic Display~
6 924 937 0 1 2
10 125
0
0 0 53872 512
6 100MEG
3 -16 45 -8
4 L160
-14 -21 14 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
4459 0 0
2
5.89979e-315 5.47595e-315
0
14 Logic Display~
6 908 937 0 1 2
10 124
0
0 0 53872 512
6 100MEG
3 -16 45 -8
3 L48
-11 -21 10 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3760 0 0
2
5.89979e-315 5.47725e-315
0
14 Logic Display~
6 892 937 0 1 2
10 123
0
0 0 53872 512
6 100MEG
3 -16 45 -8
3 L47
-11 -21 10 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
754 0 0
2
5.89979e-315 5.47854e-315
0
10 Buffer 3S~
219 419 1343 0 3 22
0 132 39 189
0
0 0 608 782
8 BUFFER3S
-27 -51 29 -43
5 U144C
-51 -5 -16 3
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
0
22

0 9 10 8 2 1 3 5 4 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 64 0
1 U
9767 0 0
2
5.89979e-315 5.47984e-315
0
8 3-In OR~
219 1199 1193 0 4 22
0 93 108 130 119
0
0 0 608 0
4 4075
-14 -24 14 -16
5 U169B
-7 -13 28 -5
0
15 DVDD=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 1 2 8 9 3 4 5 6 1
2 8 9 11 12 13 10 0 0 0
0 1 0
65 0 0 0 3 2 74 0
1 U
7978 0 0
2
5.89979e-315 5.48113e-315
0
8 3-In OR~
219 1201 1162 0 4 22
0 94 109 129 120
0
0 0 608 0
4 4075
-14 -24 14 -16
5 U169A
-7 -13 28 -5
0
15 DVDD=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 3 4 5 6 3 4 5 6 1
2 8 9 11 12 13 10 0 0 0
0 1 0
65 0 0 0 3 1 74 0
1 U
3142 0 0
2
5.89979e-315 5.48243e-315
0
8 3-In OR~
219 1202 1131 0 4 22
0 95 110 128 121
0
0 0 608 0
4 4075
-14 -24 14 -16
5 U127C
-7 -13 28 -5
0
15 DVDD=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 11 12 13 10 3 4 5 6 1
2 8 9 11 12 13 10 0 0 0
0 1 0
65 0 0 0 3 3 46 0
1 U
3284 0 0
2
5.89979e-315 5.48372e-315
0
8 3-In OR~
219 1204 1100 0 4 22
0 96 111 127 122
0
0 0 608 0
4 4075
-14 -24 14 -16
5 U127B
-7 -13 28 -5
0
15 DVDD=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 1 2 8 9 3 4 5 6 1
2 8 9 11 12 13 10 0 0 0
0 1 0
65 0 0 0 3 2 46 0
1 U
659 0 0
2
5.89979e-315 5.48502e-315
0
9 Inverter~
13 727 1424 0 2 22
0 50 51
0
0 0 608 0
6 74LS04
-21 -19 21 -11
3 z3F
-10 -3 11 5
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 13 12 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 6 68 0
1 U
3800 0 0
2
5.89979e-315 5.48631e-315
0
9 Inverter~
13 1332 1311 0 2 22
0 2 131
0
0 0 608 0
6 74LS04
-21 -19 21 -11
3 z3E
-10 -3 11 5
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 11 10 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 5 68 0
1 U
6792 0 0
2
5.89979e-315 5.48761e-315
0
12 Quad D Flop~
47 1395 1371 0 9 19
0 67 68 69 70 137 136 135 134 133
0
0 0 4704 602
4 QDFF
-14 -44 14 -36
4 U162
40 -5 68 3
0
15 DVCC=16;DGND=8;
85 %D [%16bi %8bi %1i %2i %3i %4i %9i]
+ [%16bo %1o %2o %3o %4o %9o %5o %6o %7o %8o] %M
0
11 typeDigital
5 DIP16
19

0 1 2 3 4 5 6 7 8 9
1 2 3 4 5 6 7 8 9 0
65 0 0 0 1 0 0 0
1 U
3701 0 0
2
5.89979e-315 5.4889e-315
0
13 Quad 3-State~
48 1392 1308 0 9 19
0 137 136 135 134 127 128 129 130 131
0
0 0 4704 602
8 QUAD3STA
-28 -44 28 -36
4 U165
43 -2 71 6
0
15 DVCC=16;DGND=8;
85 %D [%16bi %8bi %1i %2i %3i %4i %9i]
+ [%16bo %1o %2o %3o %4o %9o %5o %6o %7o %8o] %M
0
12 type:digital
5 DIP16
19

0 1 2 3 4 5 6 7 8 9
1 2 3 4 5 6 7 8 9 0
65 0 0 0 1 0 0 0
1 U
6316 0 0
2
5.89979e-315 5.4902e-315
0
9 2-In AND~
219 680 1910 0 3 22
0 3 102 77
0
0 0 608 0
6 74LS08
-21 -24 21 -16
5 U156D
-19 -25 16 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 67 0
1 U
8734 0 0
2
5.89979e-315 5.49149e-315
0
9 Inverter~
13 729 1910 0 2 22
0 77 138
0
0 0 608 692
6 74LS04
-21 -19 21 -11
5 U140B
-18 -20 17 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 3 4 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 2 55 0
1 U
7988 0 0
2
5.89979e-315 5.49279e-315
0
9 Inverter~
13 917 694 0 2 22
0 20 24
0
0 0 608 0
6 74LS04
-21 -19 21 -11
2 zB
-8 -6 6 2
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 3 4 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 2 66 0
1 U
3217 0 0
2
44286.3 62
0
7 Pulser~
4 671 723 0 10 12
0 616 617 18 618 0 0 5 5 6
7
0
0 0 4640 0
0
2 V5
-7 -28 7 -20
0
0
0
0
0
4 SIP2
9

0 1 2 3 4 1 2 3 4 0
0 0 0 512 1 0 0 0
1 V
3965 0 0
2
44286.3 63
0
4 4008
219 1114 557 0 14 29
0 42 47 48 49 619 620 621 11 622
140 139 118 41 623
0
0 0 4832 0
4 4008
-14 -60 14 -52
4 U153
-14 -61 14 -53
0
15 DVDD=16;DGND=8;
126 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 1 3 5 7 15 2 4 6 9
10 11 12 13 14 1 3 5 7 15
2 4 6 9 10 11 12 13 14 0
65 0 0 512 1 0 0 0
1 U
8239 0 0
2
44286.3 64
0
14 Logic Display~
6 815 486 0 1 2
10 44
0
0 0 53872 512
6 100MEG
3 -16 45 -8
3 L46
-11 -21 10 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
828 0 0
2
44286.3 65
0
10 Buffer 3S~
219 888 519 0 3 22
0 44 9 20
0
0 0 608 0
8 BUFFER3S
-27 -51 29 -43
5 U144B
-18 -20 17 -12
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
0
22

0 5 4 6 2 1 3 5 4 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 64 0
1 U
6187 0 0
2
44286.3 66
0
12 D Flip-Flop~
219 778 555 0 4 9
0 140 18 624 44
0
0 0 4704 0
3 DFF
-10 -53 11 -45
4 U147
-14 -55 14 -47
0
14 DVCC=6;DGND=5;
47 %D [%6bi %5bi %1i %2i][%6bo %1o %2o %3o %4o] %M
0
11 typeDigital
4 DIP6
9

0 1 2 3 4 1 2 3 4 0
65 0 0 512 1 0 0 0
1 U
7107 0 0
2
44286.3 67
0
14 Logic Display~
6 814 386 0 1 2
10 45
0
0 0 53872 512
6 100MEG
3 -16 45 -8
3 L43
-11 -21 10 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
6433 0 0
2
44286.3 68
0
10 Buffer 3S~
219 885 419 0 3 22
0 45 9 19
0
0 0 608 0
8 BUFFER3S
-27 -51 29 -43
5 U144A
-18 -20 17 -12
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
0
22

0 2 1 3 2 1 3 5 4 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 64 0
1 U
8559 0 0
2
44286.3 69
0
12 D Flip-Flop~
219 775 455 0 4 9
0 139 18 625 45
0
0 0 4704 0
3 DFF
-10 -53 11 -45
4 U146
-14 -55 14 -47
0
14 DVCC=6;DGND=5;
47 %D [%6bi %5bi %1i %2i][%6bo %1o %2o %3o %4o] %M
0
11 typeDigital
4 DIP6
9

0 1 2 3 4 1 2 3 4 0
65 0 0 512 1 0 0 0
1 U
3674 0 0
2
44286.3 70
0
9 Inverter~
13 339 899 0 2 22
0 50 114
0
0 0 608 0
6 74LS04
-21 -19 21 -11
5 U140C
-18 -20 17 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 5 6 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 3 55 0
1 U
5697 0 0
2
44286.3 71
0
13 Quad 3-State~
48 276 842 0 9 19
0 148 147 141 146 152 151 150 149 40
0
0 0 4704 0
8 QUAD3STA
-28 -44 28 -36
4 U163
-14 -46 14 -38
0
15 DVCC=16;DGND=8;
85 %D [%16bi %8bi %1i %2i %3i %4i %9i]
+ [%16bo %1o %2o %3o %4o %9o %5o %6o %7o %8o] %M
0
12 type:digital
5 DIP16
19

0 1 2 3 4 5 6 7 8 9
1 2 3 4 5 6 7 8 9 0
65 0 0 0 1 0 0 0
1 U
3805 0 0
2
44286.3 72
0
12 D Flip-Flop~
219 138 642 0 4 9
0 143 132 626 147
0
0 0 4704 0
3 DFF
-10 -53 11 -45
4 U161
-14 -55 14 -47
0
14 DVCC=6;DGND=5;
47 %D [%6bi %5bi %1i %2i][%6bo %1o %2o %3o %4o] %M
0
11 typeDigital
4 DIP6
9

0 1 2 3 4 1 2 3 4 0
65 0 0 512 1 0 0 0
1 U
5219 0 0
2
44286.3 73
0
10 Buffer 3S~
219 248 606 0 3 22
0 147 9 57
0
0 0 608 0
8 BUFFER3S
-27 -51 29 -43
5 U160A
-18 -20 17 -12
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
0
22

0 2 1 3 2 1 3 5 4 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 22 0
1 U
3795 0 0
2
44286.3 74
0
14 Logic Display~
6 193 573 0 1 2
10 147
0
0 0 53872 512
6 100MEG
3 -16 45 -8
4 L116
-14 -21 14 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3637 0 0
2
44286.3 75
0
14 Logic Display~
6 195 668 0 1 2
10 148
0
0 0 53872 512
6 100MEG
3 -16 45 -8
4 L115
-14 -21 14 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3226 0 0
2
44286.3 76
0
10 Buffer 3S~
219 250 701 0 3 22
0 148 9 58
0
0 0 608 0
8 BUFFER3S
-27 -51 29 -43
5 U158A
-18 -20 17 -12
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
0
22

0 2 1 3 2 1 3 5 4 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 21 0
1 U
6966 0 0
2
44286.3 77
0
12 D Flip-Flop~
219 140 737 0 4 9
0 142 132 627 148
0
0 0 4704 0
3 DFF
-10 -53 11 -45
4 U155
-14 -55 14 -47
0
14 DVCC=6;DGND=5;
47 %D [%6bi %5bi %1i %2i][%6bo %1o %2o %3o %4o] %M
0
11 typeDigital
4 DIP6
9

0 1 2 3 4 1 2 3 4 0
65 0 0 512 1 0 0 0
1 U
9796 0 0
2
44286.3 78
0
12 D Flip-Flop~
219 138 552 0 4 9
0 144 132 628 141
0
0 0 4704 0
3 DFF
-10 -53 11 -45
3 U78
-11 -55 10 -47
0
14 DVCC=6;DGND=5;
47 %D [%6bi %5bi %1i %2i][%6bo %1o %2o %3o %4o] %M
0
11 typeDigital
4 DIP6
9

0 1 2 3 4 1 2 3 4 0
65 0 0 512 1 0 0 0
1 U
5952 0 0
2
44286.3 79
0
10 Buffer 3S~
219 248 516 0 3 22
0 141 9 56
0
0 0 608 0
8 BUFFER3S
-27 -51 29 -43
5 U148D
-18 -20 17 -12
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
0
22

0 12 13 11 2 1 3 5 4 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 59 0
1 U
3649 0 0
2
44286.3 80
0
14 Logic Display~
6 193 483 0 1 2
10 141
0
0 0 53872 512
6 100MEG
3 -16 45 -8
4 L114
-14 -21 14 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3716 0 0
2
44286.3 81
0
14 Logic Display~
6 191 388 0 1 2
10 146
0
0 0 53872 512
6 100MEG
3 -16 45 -8
4 L113
-14 -21 14 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
4797 0 0
2
44286.3 82
0
10 Buffer 3S~
219 246 421 0 3 22
0 146 9 55
0
0 0 608 0
8 BUFFER3S
-27 -51 29 -43
5 U148C
-18 -20 17 -12
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
0
22

0 9 10 8 2 1 3 5 4 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 59 0
1 U
4681 0 0
2
44286.3 83
0
12 D Flip-Flop~
219 136 457 0 4 9
0 145 132 629 146
0
0 0 4704 0
3 DFF
-10 -53 11 -45
3 U77
-11 -55 10 -47
0
14 DVCC=6;DGND=5;
47 %D [%6bi %5bi %1i %2i][%6bo %1o %2o %3o %4o] %M
0
11 typeDigital
4 DIP6
9

0 1 2 3 4 1 2 3 4 0
65 0 0 512 1 0 0 0
1 U
9730 0 0
2
44286.3 84
0
4 4008
219 433 740 0 14 29
0 149 150 151 152 630 631 116 115 632
142 143 144 145 633
0
0 0 4832 0
4 4008
-14 -60 14 -52
4 U159
-14 -61 14 -53
0
15 DVDD=16;DGND=8;
126 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 1 3 5 7 15 2 4 6 9
10 11 12 13 14 1 3 5 7 15
2 4 6 9 10 11 12 13 14 0
65 0 0 512 1 0 0 0
1 U
9874 0 0
2
44286.3 85
0
10 Buffer 3S~
219 3081 1681 0 3 22
0 153 9 154
0
0 0 608 270
8 BUFFER3S
-27 -51 29 -43
5 U148B
13 -5 48 3
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
0
22

0 5 4 6 2 1 3 5 4 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 59 0
1 U
364 0 0
2
44286.3 86
0
9 2-In AND~
219 3060 1481 0 3 22
0 90 157 158
0
0 0 608 180
6 74LS08
-21 -24 21 -16
5 U152D
-19 -2 16 6
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 63 0
1 U
3656 0 0
2
44286.3 87
0
9 2-In AND~
219 2732 1485 0 3 22
0 90 159 160
0
0 0 608 180
6 74LS08
-21 -24 21 -16
5 U152C
-19 -2 16 6
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 63 0
1 U
3131 0 0
2
44286.3 88
0
9 2-In AND~
219 2444 1480 0 3 22
0 90 161 162
0
0 0 608 180
6 74LS08
-21 -24 21 -16
5 U152B
-19 -2 16 6
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 63 0
1 U
6772 0 0
2
44286.3 89
0
9 2-In AND~
219 2155 1484 0 3 22
0 90 163 164
0
0 0 608 180
6 74LS08
-21 -24 21 -16
5 U152A
-19 -2 16 6
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 63 0
1 U
9557 0 0
2
44286.3 90
0
9 2-In AND~
219 3064 1250 0 3 22
0 90 165 166
0
0 0 608 180
6 74LS08
-21 -24 21 -16
5 U151D
-19 -2 16 6
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 62 0
1 U
5789 0 0
2
44286.3 91
0
9 2-In AND~
219 2741 1249 0 3 22
0 90 167 168
0
0 0 608 180
6 74LS08
-21 -24 21 -16
5 U151C
-19 -2 16 6
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 62 0
1 U
7328 0 0
2
44286.3 92
0
9 2-In AND~
219 2455 1250 0 3 22
0 90 169 170
0
0 0 608 180
6 74LS08
-21 -24 21 -16
5 U151B
-19 -2 16 6
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 62 0
1 U
4799 0 0
2
44286.3 93
0
9 2-In AND~
219 2165 1254 0 3 22
0 90 171 172
0
0 0 608 180
6 74LS08
-21 -24 21 -16
5 U151A
-19 -2 16 6
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 62 0
1 U
9196 0 0
2
44286.3 94
0
9 2-In AND~
219 3053 1033 0 3 22
0 90 173 174
0
0 0 608 180
6 74LS08
-21 -24 21 -16
5 U150D
-19 -2 16 6
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 61 0
1 U
3857 0 0
2
44286.3 95
0
9 2-In AND~
219 2737 1037 0 3 22
0 90 175 176
0
0 0 608 180
6 74LS08
-21 -24 21 -16
5 U150C
-19 -2 16 6
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 61 0
1 U
7125 0 0
2
44286.3 96
0
9 2-In AND~
219 2453 1029 0 3 22
0 90 177 178
0
0 0 608 180
6 74LS08
-21 -24 21 -16
5 U150B
-19 -2 16 6
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 61 0
1 U
3641 0 0
2
44286.3 97
0
9 2-In AND~
219 2167 1037 0 3 22
0 90 179 180
0
0 0 608 180
6 74LS08
-21 -24 21 -16
5 U150A
-19 -2 16 6
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 61 0
1 U
9821 0 0
2
44286.3 98
0
9 2-In AND~
219 3054 811 0 3 22
0 90 181 182
0
0 0 608 180
6 74LS08
-21 -24 21 -16
5 U149D
-19 -2 16 6
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 60 0
1 U
3187 0 0
2
44286.3 99
0
9 2-In AND~
219 2743 812 0 3 22
0 90 183 184
0
0 0 608 180
6 74LS08
-21 -24 21 -16
5 U149C
-19 -2 16 6
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 60 0
1 U
762 0 0
2
44286.3 100
0
9 2-In AND~
219 2461 812 0 3 22
0 90 186 187
0
0 0 608 180
6 74LS08
-21 -24 21 -16
5 U149B
-19 -2 16 6
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 60 0
1 U
39 0 0
2
44286.3 101
0
9 2-In AND~
219 2172 814 0 3 22
0 90 185 188
0
0 0 608 180
6 74LS08
-21 -24 21 -16
5 U149A
-19 -2 16 6
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 60 0
1 U
9450 0 0
2
44286.3 102
0
4 4008
219 1132 1343 0 14 29
0 97 98 99 100 634 635 636 117 637
104 105 106 107 638
0
0 0 4832 0
4 4008
-14 -60 14 -52
4 U145
-14 -61 14 -53
0
15 DVDD=16;DGND=8;
126 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 1 3 5 7 15 2 4 6 9
10 11 12 13 14 1 3 5 7 15
2 4 6 9 10 11 12 13 14 0
65 0 0 512 1 0 0 0
1 U
3236 0 0
2
44286.3 103
0
13 Quad 3-State~
48 726 1820 0 9 19
0 67 68 69 70 193 192 191 190 138
0
0 0 4704 270
8 QUAD3STA
-28 -44 28 -36
4 U142
39 -1 67 7
0
15 DVCC=16;DGND=8;
85 %D [%16bi %8bi %1i %2i %3i %4i %9i]
+ [%16bo %1o %2o %3o %4o %9o %5o %6o %7o %8o] %M
0
12 type:digital
5 DIP16
19

0 1 2 3 4 5 6 7 8 9
1 2 3 4 5 6 7 8 9 0
65 0 0 0 1 0 0 0
1 U
3321 0 0
2
5.89979e-315 5.49408e-315
0
8 2-In OR~
219 1253 2904 0 3 22
0 200 198 199
0
0 0 608 90
6 74LS32
-21 -24 21 -16
4 U94D
29 -3 57 5
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 51 0
1 U
8879 0 0
2
5.89979e-315 5.49538e-315
0
13 Quad 3-State~
48 1894 3190 0 9 19
0 227 228 229 230 202 203 204 205 231
0
0 0 4704 692
8 QUAD3STA
-28 -44 28 -36
4 U138
-14 46 14 54
0
15 DVCC=16;DGND=8;
85 %D [%16bi %8bi %1i %2i %3i %4i %9i]
+ [%16bo %1o %2o %3o %4o %9o %5o %6o %7o %8o] %M
0
12 type:digital
5 DIP16
19

0 4 5 12 13 2 7 10 15 9
4 5 12 13 2 7 10 15 9 0
65 0 0 0 1 0 0 0
1 U
5433 0 0
2
44286.3 104
0
9 Inverter~
13 1871 3139 0 2 22
0 198 231
0
0 0 608 692
6 74LS04
-21 -19 21 -11
5 U132F
-18 -20 17 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 13 12 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 6 49 0
1 U
3679 0 0
2
44286.3 105
0
14 Logic Display~
6 1937 3161 0 1 2
10 205
0
0 0 53872 512
6 100MEG
3 -16 45 -8
3 L16
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
9342 0 0
2
44286.3 106
0
14 Logic Display~
6 1950 3161 0 1 2
10 204
0
0 0 53872 512
6 100MEG
3 -16 45 -8
3 L15
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3623 0 0
2
44286.3 107
0
14 Logic Display~
6 1963 3162 0 1 2
10 203
0
0 0 53872 512
6 100MEG
3 -16 45 -8
3 L14
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3722 0 0
2
44286.3 108
0
14 Logic Display~
6 1976 3162 0 1 2
10 202
0
0 0 53872 512
6 100MEG
3 -16 45 -8
3 L13
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
8993 0 0
2
44286.3 109
0
5 4030~
219 1696 3164 0 3 22
0 225 221 230
0
0 0 608 0
4 4030
-7 -24 21 -16
5 U137C
-6 -15 29 -7
0
15 DVDD=14;DGND=7;
49 %D [%14bi %7bi %1i %2i]
+ [%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 8 9 10 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 3 54 0
1 U
3723 0 0
2
44286.3 110
0
5 4030~
219 1696 3197 0 3 22
0 224 220 229
0
0 0 608 0
4 4030
-7 -24 21 -16
5 U137B
-4 -16 31 -8
0
15 DVDD=14;DGND=7;
49 %D [%14bi %7bi %1i %2i]
+ [%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 5 6 4 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 2 54 0
1 U
6244 0 0
2
44286.3 111
0
5 4030~
219 1696 3231 0 3 22
0 223 219 228
0
0 0 608 0
4 4030
-7 -24 21 -16
5 U137A
-3 -13 32 -5
0
15 DVDD=14;DGND=7;
49 %D [%14bi %7bi %1i %2i]
+ [%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 1 54 0
1 U
6421 0 0
2
44286.3 112
0
5 4030~
219 1695 3266 0 3 22
0 222 218 227
0
0 0 608 0
4 4030
-7 -24 21 -16
5 U117A
-2 -11 33 -3
0
15 DVDD=14;DGND=7;
49 %D [%14bi %7bi %1i %2i]
+ [%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 1 52 0
1 U
7743 0 0
2
44286.3 113
0
5 4030~
219 1695 3081 0 3 22
0 16 222 232
0
0 0 608 0
4 4030
-7 -24 21 -16
5 U136D
-2 -11 33 -3
0
15 DVDD=14;DGND=7;
49 %D [%14bi %7bi %1i %2i]
+ [%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 4 53 0
1 U
9840 0 0
2
44286.3 114
0
5 4030~
219 1696 3046 0 3 22
0 15 223 233
0
0 0 608 0
4 4030
-7 -24 21 -16
5 U136C
-3 -13 32 -5
0
15 DVDD=14;DGND=7;
49 %D [%14bi %7bi %1i %2i]
+ [%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 8 9 10 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 3 53 0
1 U
6910 0 0
2
44286.3 115
0
5 4030~
219 1696 3012 0 3 22
0 14 224 234
0
0 0 608 0
4 4030
-7 -24 21 -16
5 U136B
-4 -16 31 -8
0
15 DVDD=14;DGND=7;
49 %D [%14bi %7bi %1i %2i]
+ [%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 5 6 4 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 2 53 0
1 U
449 0 0
2
44286.3 116
0
5 4030~
219 1696 2979 0 3 22
0 13 225 235
0
0 0 608 0
4 4030
-7 -24 21 -16
5 U136A
-6 -15 29 -7
0
15 DVDD=14;DGND=7;
49 %D [%14bi %7bi %1i %2i]
+ [%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 1 53 0
1 U
8761 0 0
2
44286.3 117
0
14 Logic Display~
6 1976 2977 0 1 2
10 206
0
0 0 53872 512
6 100MEG
3 -16 45 -8
3 L12
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
6748 0 0
2
44286.3 118
0
14 Logic Display~
6 1963 2977 0 1 2
10 207
0
0 0 53872 512
6 100MEG
3 -16 45 -8
3 L11
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
7393 0 0
2
44286.3 119
0
14 Logic Display~
6 1950 2976 0 1 2
10 208
0
0 0 53872 512
6 100MEG
3 -16 45 -8
3 L10
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
7699 0 0
2
44286.3 120
0
14 Logic Display~
6 1937 2976 0 1 2
10 209
0
0 0 53872 512
6 100MEG
3 -16 45 -8
2 L9
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
6638 0 0
2
44286.3 121
0
9 Inverter~
13 1871 2954 0 2 22
0 200 236
0
0 0 608 692
6 74LS04
-21 -19 21 -11
5 U132E
-18 -20 17 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 11 10 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 5 49 0
1 U
4595 0 0
2
44286.3 122
0
13 Quad 3-State~
48 1894 3005 0 9 19
0 232 233 234 235 206 207 208 209 236
0
0 0 4704 692
8 QUAD3STA
-28 -44 28 -36
4 U135
-14 46 14 54
0
15 DVCC=16;DGND=8;
85 %D [%16bi %8bi %1i %2i %3i %4i %9i]
+ [%16bo %1o %2o %3o %4o %9o %5o %6o %7o %8o] %M
0
12 type:digital
5 DIP16
19

0 4 5 12 13 2 7 10 15 9
4 5 12 13 2 7 10 15 9 0
65 0 0 0 1 0 0 0
1 U
9395 0 0
2
44286.3 123
0
8 2-In OR~
219 1694 2782 0 3 22
0 225 221 240
0
0 0 608 0
6 74LS32
-21 -24 21 -16
4 U94C
-3 -14 25 -6
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 9 10 8 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 51 0
1 U
3303 0 0
2
44286.3 124
0
8 2-In OR~
219 1694 2815 0 3 22
0 224 220 239
0
0 0 608 0
6 74LS32
-21 -24 21 -16
4 U94B
0 -14 28 -6
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 51 0
1 U
4498 0 0
2
44286.3 125
0
8 2-In OR~
219 1694 2850 0 3 22
0 223 219 238
0
0 0 608 0
6 74LS32
-21 -24 21 -16
4 U94A
-3 -12 25 -4
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 51 0
1 U
9728 0 0
2
44286.3 126
0
8 2-In OR~
219 1694 2884 0 3 22
0 222 218 237
0
0 0 608 0
6 74LS32
-21 -24 21 -16
4 U93A
-3 -12 25 -4
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 41 0
1 U
3789 0 0
2
44286.3 127
0
13 Quad 3-State~
48 1891 2808 0 9 19
0 237 238 239 240 210 211 212 213 241
0
0 0 4704 692
8 QUAD3STA
-28 -44 28 -36
3 U35
-11 46 10 54
0
15 DVCC=16;DGND=8;
85 %D [%16bi %8bi %1i %2i %3i %4i %9i]
+ [%16bo %1o %2o %3o %4o %9o %5o %6o %7o %8o] %M
0
12 type:digital
5 DIP16
19

0 4 5 12 13 2 7 10 15 9
4 5 12 13 2 7 10 15 9 0
65 0 0 0 1 0 0 0
1 U
3978 0 0
2
44286.3 128
0
9 Inverter~
13 1868 2757 0 2 22
0 201 241
0
0 0 608 692
6 74LS04
-21 -19 21 -11
5 U132D
-18 -20 17 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 9 8 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 4 49 0
1 U
3494 0 0
2
44286.3 129
0
14 Logic Display~
6 1934 2779 0 1 2
10 213
0
0 0 53872 512
6 100MEG
3 -16 45 -8
2 L8
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3507 0 0
2
44286.3 130
0
14 Logic Display~
6 1947 2779 0 1 2
10 212
0
0 0 53872 512
6 100MEG
3 -16 45 -8
2 L7
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
5151 0 0
2
44286.3 131
0
14 Logic Display~
6 1960 2780 0 1 2
10 211
0
0 0 53872 512
6 100MEG
3 -16 45 -8
2 L6
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3701 0 0
2
44286.3 132
0
14 Logic Display~
6 1973 2780 0 1 2
10 210
0
0 0 53872 512
6 100MEG
3 -16 45 -8
2 L5
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
8585 0 0
2
44286.3 133
0
14 Logic Display~
6 1972 2599 0 1 2
10 214
0
0 0 53872 512
6 100MEG
3 -16 45 -8
2 L4
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
8809 0 0
2
44286.3 134
0
14 Logic Display~
6 1959 2599 0 1 2
10 215
0
0 0 53872 512
6 100MEG
3 -16 45 -8
2 L3
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
5993 0 0
2
44286.3 135
0
14 Logic Display~
6 1946 2598 0 1 2
10 216
0
0 0 53872 512
6 100MEG
3 -16 45 -8
2 L2
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
8654 0 0
2
44286.3 136
0
14 Logic Display~
6 1933 2598 0 1 2
10 217
0
0 0 53872 512
6 100MEG
3 -16 45 -8
2 L1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
7223 0 0
2
44286.3 137
0
9 Inverter~
13 1867 2576 0 2 22
0 226 246
0
0 0 608 692
6 74LS04
-21 -19 21 -11
5 U132C
-18 -20 17 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 5 6 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 3 49 0
1 U
3641 0 0
2
44286.3 138
0
13 Quad 3-State~
48 1890 2627 0 9 19
0 242 243 244 245 214 215 216 217 246
0
0 0 4704 692
8 QUAD3STA
-28 -44 28 -36
3 U10
-11 46 10 54
0
15 DVCC=16;DGND=8;
85 %D [%16bi %8bi %1i %2i %3i %4i %9i]
+ [%16bo %1o %2o %3o %4o %9o %5o %6o %7o %8o] %M
0
12 type:digital
5 DIP16
19

0 4 5 12 13 2 7 10 15 9
4 5 12 13 2 7 10 15 9 0
65 0 0 0 1 0 0 0
1 U
3104 0 0
2
44286.3 139
0
14 Logic Display~
6 2503 2718 0 1 2
10 250
0
0 0 53872 512
6 100MEG
3 -16 45 -8
4 L159
-14 -21 14 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3296 0 0
2
44286.3 140
0
14 Logic Display~
6 2516 2718 0 1 2
10 249
0
0 0 53872 512
6 100MEG
3 -16 45 -8
4 L158
-14 -21 14 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
8534 0 0
2
44286.3 141
0
14 Logic Display~
6 2529 2719 0 1 2
10 248
0
0 0 53872 512
6 100MEG
3 -16 45 -8
4 L157
-14 -21 14 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
949 0 0
2
44286.3 142
0
14 Logic Display~
6 2542 2719 0 1 2
10 247
0
0 0 53872 512
6 100MEG
3 -16 45 -8
4 L156
-14 -21 14 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3371 0 0
2
44286.3 143
0
14 Logic Display~
6 2500 2540 0 1 2
10 254
0
0 0 53872 512
6 100MEG
3 -16 45 -8
4 L155
-14 -21 14 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
7311 0 0
2
44286.3 144
0
14 Logic Display~
6 2513 2540 0 1 2
10 253
0
0 0 53872 512
6 100MEG
3 -16 45 -8
4 L154
-14 -21 14 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3409 0 0
2
44286.3 145
0
14 Logic Display~
6 2526 2541 0 1 2
10 252
0
0 0 53872 512
6 100MEG
3 -16 45 -8
4 L153
-14 -21 14 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3526 0 0
2
44286.3 146
0
14 Logic Display~
6 2539 2541 0 1 2
10 251
0
0 0 53872 512
6 100MEG
3 -16 45 -8
4 L152
-14 -21 14 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
4129 0 0
2
44286.3 147
0
14 Logic Display~
6 2538 2345 0 1 2
10 256
0
0 0 53872 512
6 100MEG
3 -16 45 -8
4 L148
-14 -21 14 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
6278 0 0
2
44286.3 148
0
14 Logic Display~
6 2525 2345 0 1 2
10 257
0
0 0 53872 512
6 100MEG
3 -16 45 -8
4 L149
-14 -21 14 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3482 0 0
2
44286.3 149
0
14 Logic Display~
6 2512 2344 0 1 2
10 258
0
0 0 53872 512
6 100MEG
3 -16 45 -8
4 L150
-14 -21 14 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
8323 0 0
2
44286.3 150
0
14 Logic Display~
6 2499 2344 0 1 2
10 259
0
0 0 53872 512
6 100MEG
3 -16 45 -8
4 L151
-14 -21 14 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3984 0 0
2
44286.3 151
0
13 Quad 3-State~
48 2459 2747 0 9 19
0 261 262 263 264 247 248 249 250 265
0
0 0 4704 692
8 QUAD3STA
-28 -44 28 -36
4 U134
-14 46 14 54
0
15 DVCC=16;DGND=8;
85 %D [%16bi %8bi %1i %2i %3i %4i %9i]
+ [%16bo %1o %2o %3o %4o %9o %5o %6o %7o %8o] %M
0
12 type:digital
5 DIP16
19

0 4 5 12 13 2 7 10 15 9
4 5 12 13 2 7 10 15 9 0
65 0 0 0 1 0 0 0
1 U
7622 0 0
2
44286.3 152
0
9 2-In AND~
219 2272 2721 0 3 22
0 221 13 264
0
0 0 608 0
6 74LS08
-21 -24 21 -16
5 U133D
-13 -8 22 0
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 50 0
1 U
816 0 0
2
44286.3 153
0
9 2-In AND~
219 2272 2755 0 3 22
0 220 14 263
0
0 0 608 0
6 74LS08
-21 -24 21 -16
5 U133C
-17 -11 18 -3
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 50 0
1 U
4656 0 0
2
44286.3 154
0
9 2-In AND~
219 2274 2822 0 3 22
0 218 16 261
0
0 0 608 0
6 74LS08
-21 -24 21 -16
5 U133B
-13 -12 22 -4
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 50 0
1 U
6356 0 0
2
44286.3 155
0
9 2-In AND~
219 2273 2788 0 3 22
0 219 15 262
0
0 0 608 0
6 74LS08
-21 -24 21 -16
5 U133A
-13 -11 22 -3
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 50 0
1 U
7479 0 0
2
44286.3 156
0
9 Inverter~
13 2436 2696 0 2 22
0 255 265
0
0 0 608 692
6 74LS04
-21 -19 21 -11
5 U132B
-18 -20 17 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 3 4 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 2 49 0
1 U
5690 0 0
2
44286.3 157
0
13 Quad 3-State~
48 2456 2569 0 9 19
0 266 267 268 269 251 252 253 254 270
0
0 0 4704 692
8 QUAD3STA
-28 -44 28 -36
3 U97
-11 46 10 54
0
15 DVCC=16;DGND=8;
85 %D [%16bi %8bi %1i %2i %3i %4i %9i]
+ [%16bo %1o %2o %3o %4o %9o %5o %6o %7o %8o] %M
0
12 type:digital
5 DIP16
19

0 4 5 12 13 2 7 10 15 9
4 5 12 13 2 7 10 15 9 0
65 0 0 0 1 0 0 0
1 U
5617 0 0
2
44286.3 158
0
9 2-In AND~
219 2269 2543 0 3 22
0 225 221 269
0
0 0 608 0
6 74LS08
-21 -24 21 -16
5 U129C
-15 -10 20 -2
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 48 0
1 U
3903 0 0
2
44286.3 159
0
9 2-In AND~
219 2270 2577 0 3 22
0 224 220 268
0
0 0 608 0
6 74LS08
-21 -24 21 -16
5 U129D
-16 -13 19 -5
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 48 0
1 U
4452 0 0
2
44286.3 160
0
9 2-In AND~
219 2271 2644 0 3 22
0 222 218 266
0
0 0 608 0
6 74LS08
-21 -24 21 -16
5 U130A
-16 -12 19 -4
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 34 0
1 U
6282 0 0
2
44286.3 161
0
9 2-In AND~
219 2270 2610 0 3 22
0 223 219 267
0
0 0 608 0
6 74LS08
-21 -24 21 -16
5 U131A
-17 -13 18 -5
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 35 0
1 U
7187 0 0
2
44286.3 162
0
9 Inverter~
13 2433 2518 0 2 22
0 260 270
0
0 0 608 692
6 74LS04
-21 -19 21 -11
5 U132A
-18 -20 17 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 1 49 0
1 U
6866 0 0
2
44286.3 163
0
8 2-In OR~
219 1693 2703 0 3 22
0 16 222 242
0
0 0 608 0
6 74LS32
-21 -24 21 -16
4 U99C
-3 -12 25 -4
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 9 10 8 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 37 0
1 U
7670 0 0
2
44286.3 164
0
8 2-In OR~
219 1693 2669 0 3 22
0 15 223 243
0
0 0 608 0
6 74LS32
-21 -24 21 -16
4 U99B
-3 -12 25 -4
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 37 0
1 U
951 0 0
2
44286.3 165
0
8 2-In OR~
219 1693 2634 0 3 22
0 14 224 244
0
0 0 608 0
6 74LS32
-21 -24 21 -16
4 U99A
0 -14 28 -6
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 37 0
1 U
9536 0 0
2
44286.3 166
0
8 2-In OR~
219 1693 2601 0 3 22
0 13 225 245
0
0 0 608 0
6 74LS32
-21 -24 21 -16
4 U86D
-3 -14 25 -6
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 30 0
1 U
5495 0 0
2
44286.3 167
0
9 Inverter~
13 2433 2325 0 2 22
0 275 276
0
0 0 608 692
6 74LS04
-21 -19 21 -11
5 U124F
-18 -20 17 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 13 12 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 6 44 0
1 U
8152 0 0
2
44286.3 168
0
13 Quad 3-State~
48 2454 2373 0 9 19
0 271 272 273 274 256 257 258 259 276
0
0 0 4704 692
8 QUAD3STA
-28 -44 28 -36
3 U96
-11 46 10 54
0
15 DVCC=16;DGND=8;
85 %D [%16bi %8bi %1i %2i %3i %4i %9i]
+ [%16bo %1o %2o %3o %4o %9o %5o %6o %7o %8o] %M
0
12 type:digital
5 DIP16
19

0 4 5 12 13 2 7 10 15 9
4 5 12 13 2 7 10 15 9 0
65 0 0 0 1 0 0 0
1 U
6223 0 0
2
44286.3 169
0
9 2-In AND~
219 2267 2347 0 3 22
0 13 225 274
0
0 0 608 0
6 74LS08
-21 -24 21 -16
3 U6B
-16 -9 5 -1
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 5 0
1 U
5441 0 0
2
44286.3 170
0
9 2-In AND~
219 2268 2381 0 3 22
0 14 224 273
0
0 0 608 0
6 74LS08
-21 -24 21 -16
4 U98B
-19 -9 9 -1
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 36 0
1 U
3189 0 0
2
44286.3 171
0
9 2-In AND~
219 2269 2448 0 3 22
0 16 222 271
0
0 0 608 0
6 74LS08
-21 -24 21 -16
4 U98C
-19 -9 9 -1
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 36 0
1 U
8460 0 0
2
44286.3 172
0
9 2-In AND~
219 2268 2414 0 3 22
0 15 223 272
0
0 0 608 0
6 74LS08
-21 -24 21 -16
4 U98D
-19 -9 9 -1
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 36 0
1 U
5179 0 0
2
44286.3 173
0
7 Pulser~
4 2937 2237 0 10 12
0 639 640 277 641 0 0 5 5 6
7
0
0 0 4640 0
0
3 V33
-10 -28 11 -20
0
0
0
0
0
4 SIP2
9

0 1 2 3 4 1 2 3 4 0
0 0 0 512 1 0 0 0
1 V
3593 0 0
2
44286.3 174
0
8 2-In OR~
219 2053 2109 0 3 22
0 339 338 329
0
0 0 608 0
6 74LS32
-21 -24 21 -16
5 U126D
-9 -9 26 -1
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 45 0
1 U
3928 0 0
2
44286.3 175
0
8 2-In OR~
219 2055 1966 0 3 22
0 340 339 330
0
0 0 608 0
6 74LS32
-21 -24 21 -16
5 U126C
-9 -9 26 -1
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 9 10 8 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 45 0
1 U
363 0 0
2
44286.3 176
0
8 2-In OR~
219 2054 1800 0 3 22
0 340 338 328
0
0 0 608 0
6 74LS32
-21 -24 21 -16
5 U126B
-9 -9 26 -1
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 45 0
1 U
8132 0 0
2
44286.3 177
0
9 Inverter~
13 2556 2142 0 2 22
0 294 295
0
0 0 608 602
6 74LS04
-21 -19 21 -11
5 U124E
-8 1 27 9
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 11 10 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 5 44 0
1 U
65 0 0
2
44286.3 178
0
9 Inverter~
13 2551 1970 0 2 22
0 296 297
0
0 0 608 602
6 74LS04
-21 -19 21 -11
5 U124D
-16 1 19 9
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 9 8 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 4 44 0
1 U
6609 0 0
2
44286.3 179
0
9 Inverter~
13 2567 1821 0 2 22
0 303 304
0
0 0 608 692
6 74LS04
-21 -19 21 -11
5 U124C
-18 -20 17 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 5 6 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 3 44 0
1 U
8995 0 0
2
44286.3 180
0
10 Buffer 3S~
219 2559 2117 0 3 22
0 300 295 298
0
0 0 608 0
8 BUFFER3S
-27 -51 29 -43
5 U128C
-18 -20 17 -12
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
0
22

0 9 10 8 2 1 3 5 4 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 47 0
1 U
3918 0 0
2
44286.3 181
0
10 Buffer 3S~
219 2554 1946 0 3 22
0 301 297 299
0
0 0 608 0
8 BUFFER3S
-27 -51 29 -43
5 U128B
-18 -20 17 -12
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
0
22

0 5 4 6 2 1 3 5 4 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 47 0
1 U
7519 0 0
2
44286.3 182
0
10 Buffer 3S~
219 2589 1787 0 3 22
0 302 304 305
0
0 0 608 0
8 BUFFER3S
-27 -51 29 -43
5 U128A
-18 -20 17 -12
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
0
22

0 2 1 3 2 1 3 5 4 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 47 0
1 U
377 0 0
2
44286.3 183
0
8 3-In OR~
219 2633 1812 0 4 22
0 305 299 298 306
0
0 0 608 0
4 4075
-14 -24 14 -16
5 U127A
-10 -25 25 -17
0
15 DVDD=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 3 4 5 6 3 4 5 6 1
2 8 9 11 12 13 10 0 0 0
0 1 0
65 0 0 0 3 1 46 0
1 U
8816 0 0
2
44286.3 184
0
14 Logic Display~
6 2921 2002 0 1 2
10 306
0
0 0 53872 512
6 100MEG
3 -16 45 -8
4 Cout
-14 -21 14 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3877 0 0
2
44286.3 185
0
8 2-In OR~
219 2821 2352 0 3 22
0 319 318 315
0
0 0 608 0
6 74LS32
-21 -24 21 -16
5 U126A
-9 -9 26 -1
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 45 0
1 U
926 0 0
2
44286.3 186
0
8 2-In OR~
219 2747 2352 0 3 22
0 209 205 318
0
0 0 608 0
6 74LS32
-21 -24 21 -16
5 U120D
-9 -9 26 -1
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 43 0
1 U
7262 0 0
2
44286.3 187
0
9 Inverter~
13 2805 2312 0 2 22
0 320 319
0
0 0 608 270
6 74LS04
-21 -19 21 -11
5 U124B
-15 -15 20 -7
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 3 4 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 2 44 0
1 U
5267 0 0
2
44286.3 188
0
9 8-In NOR~
219 2749 2296 0 9 19
0 213 217 250 254 259 289 290 307 320
0
0 0 608 692
4 4078
-7 -24 21 -16
4 U125
-5 -33 23 -25
0
15 DVDD=14;DGND=7;
97 %D [%14bi %7bi %1i %2i %3i %4i %5i %6i %7i %8i]
+ [%14bo %1o %2o %3o %4o %5o %6o %7o %8o %9o] %M
0
12 type:digital
5 DIP14
19

0 2 3 4 5 9 10 11 12 13
2 3 4 5 9 10 11 12 13 0
65 0 0 0 1 0 0 0
1 U
8838 0 0
2
44286.3 189
0
8 2-In OR~
219 2814 2226 0 3 22
0 322 321 316
0
0 0 608 0
6 74LS32
-21 -24 21 -16
5 U120C
-9 -9 26 -1
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 9 10 8 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 43 0
1 U
7159 0 0
2
44286.3 190
0
8 2-In OR~
219 2747 2229 0 3 22
0 208 204 321
0
0 0 608 0
6 74LS32
-21 -24 21 -16
5 U120B
-9 -9 26 -1
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 43 0
1 U
5812 0 0
2
44286.3 191
0
9 Inverter~
13 2796 2190 0 2 22
0 323 322
0
0 0 608 270
6 74LS04
-21 -19 21 -11
5 U124A
-15 -15 20 -7
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 1 44 0
1 U
331 0 0
2
44286.3 192
0
9 8-In NOR~
219 2750 2174 0 9 19
0 212 216 249 253 258 288 291 308 323
0
0 0 608 692
4 4078
-7 -24 21 -16
4 U123
-10 -27 18 -19
0
15 DVDD=14;DGND=7;
97 %D [%14bi %7bi %1i %2i %3i %4i %5i %6i %7i %8i]
+ [%14bo %1o %2o %3o %4o %5o %6o %7o %8o %9o] %M
0
12 type:digital
5 DIP14
19

0 2 3 4 5 9 10 11 12 13
2 3 4 5 9 10 11 12 13 0
65 0 0 0 1 0 0 0
1 U
9604 0 0
2
44286.3 193
0
8 2-In OR~
219 2810 2102 0 3 22
0 325 324 317
0
0 0 608 0
6 74LS32
-21 -24 21 -16
5 U120A
-9 -9 26 -1
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 43 0
1 U
7518 0 0
2
44286.3 194
0
8 2-In OR~
219 2748 2107 0 3 22
0 207 203 324
0
0 0 608 0
6 74LS32
-21 -24 21 -16
5 U111D
-9 -9 26 -1
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 40 0
1 U
4832 0 0
2
44286.3 195
0
9 Inverter~
13 2790 2068 0 2 22
0 326 325
0
0 0 608 270
6 74LS04
-21 -19 21 -11
5 U110F
-15 -15 20 -7
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 13 12 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 6 39 0
1 U
6798 0 0
2
44286.3 196
0
9 8-In NOR~
219 2751 2049 0 9 19
0 211 215 248 252 257 287 292 309 326
0
0 0 608 692
4 4078
-7 -24 21 -16
4 U115
-6 -30 22 -22
0
15 DVDD=14;DGND=7;
97 %D [%14bi %7bi %1i %2i %3i %4i %5i %6i %7i %8i]
+ [%14bo %1o %2o %3o %4o %5o %6o %7o %8o %9o] %M
0
12 type:digital
5 DIP14
19

0 2 3 4 5 9 10 11 12 13
2 3 4 5 9 10 11 12 13 0
65 0 0 0 1 0 0 0
1 U
3336 0 0
2
44286.3 197
0
13 Quad 3-State~
48 2538 2195 0 9 19
0 281 280 279 278 286 287 288 289 294
0
0 0 4704 692
8 QUAD3STA
-28 -44 28 -36
4 U122
-14 46 14 54
0
15 DVCC=16;DGND=8;
85 %D [%16bi %8bi %1i %2i %3i %4i %9i]
+ [%16bo %1o %2o %3o %4o %9o %5o %6o %7o %8o] %M
0
12 type:digital
5 DIP16
19

0 4 5 12 13 2 7 10 15 9
4 5 12 13 2 7 10 15 9 0
65 0 0 0 1 0 0 0
1 U
8370 0 0
2
44286.3 198
0
13 Quad 3-State~
48 2539 2038 0 9 19
0 285 284 283 282 293 292 291 290 296
0
0 0 4704 692
8 QUAD3STA
-28 -44 28 -36
4 U121
-14 46 14 54
0
15 DVCC=16;DGND=8;
85 %D [%16bi %8bi %1i %2i %3i %4i %9i]
+ [%16bo %1o %2o %3o %4o %9o %5o %6o %7o %8o] %M
0
12 type:digital
5 DIP16
19

0 4 5 12 13 2 7 10 15 9
4 5 12 13 2 7 10 15 9 0
65 0 0 0 1 0 0 0
1 U
3910 0 0
2
44286.3 199
0
13 Quad 3-State~
48 2540 1863 0 9 19
0 314 313 312 311 310 309 308 307 303
0
0 0 4704 692
8 QUAD3STA
-28 -44 28 -36
4 U112
-14 46 14 54
0
15 DVCC=16;DGND=8;
85 %D [%16bi %8bi %1i %2i %3i %4i %9i]
+ [%16bo %1o %2o %3o %4o %9o %5o %6o %7o %8o] %M
0
12 type:digital
5 DIP16
19

0 4 5 12 13 2 7 10 15 9
4 5 12 13 2 7 10 15 9 0
65 0 0 0 1 0 0 0
1 U
316 0 0
2
44286.3 200
0
9 8-In NOR~
219 2752 1929 0 9 19
0 210 214 247 251 256 286 293 310 333
0
0 0 608 692
4 4078
-7 -24 21 -16
4 U119
-5 -27 23 -19
0
15 DVDD=14;DGND=7;
97 %D [%14bi %7bi %1i %2i %3i %4i %5i %6i %7i %8i]
+ [%14bo %1o %2o %3o %4o %5o %6o %7o %8o %9o] %M
0
12 type:digital
5 DIP14
19

0 2 3 4 5 9 10 11 12 13
2 3 4 5 9 10 11 12 13 0
65 0 0 0 1 0 0 0
1 U
536 0 0
2
5.89979e-315 5.49667e-315
0
9 Inverter~
13 2796 1948 0 2 22
0 333 332
0
0 0 608 270
6 74LS04
-21 -19 21 -11
5 U110E
-15 -15 20 -7
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 11 10 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 5 39 0
1 U
4460 0 0
2
5.89979e-315 5.49797e-315
0
8 2-In OR~
219 2750 1981 0 3 22
0 206 202 331
0
0 0 608 0
6 74LS32
-21 -24 21 -16
5 U111B
-9 -9 26 -1
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 40 0
1 U
3260 0 0
2
5.89979e-315 5.49926e-315
0
8 2-In OR~
219 2817 1976 0 3 22
0 332 331 327
0
0 0 608 0
6 74LS32
-21 -24 21 -16
5 U111C
-9 -9 26 -1
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 9 10 8 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 40 0
1 U
5156 0 0
2
5.89979e-315 5.50056e-315
0
14 Logic Display~
6 2993 2002 0 1 2
10 337
0
0 0 53872 512
6 100MEG
3 -16 45 -8
4 L125
-14 -21 14 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3133 0 0
2
5.89979e-315 5.50185e-315
0
14 Logic Display~
6 2980 2002 0 1 2
10 336
0
0 0 53872 512
6 100MEG
3 -16 45 -8
4 L126
-14 -21 14 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
5523 0 0
2
5.89979e-315 5.50315e-315
0
14 Logic Display~
6 2967 2002 0 1 2
10 335
0
0 0 53872 512
6 100MEG
3 -16 45 -8
4 L127
-14 -21 14 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3746 0 0
2
5.89979e-315 5.50444e-315
0
14 Logic Display~
6 2954 2002 0 1 2
10 334
0
0 0 53872 512
6 100MEG
3 -16 45 -8
4 L128
-14 -21 14 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
5668 0 0
2
5.89979e-315 5.50574e-315
0
12 Quad D Flop~
47 2884 2071 0 9 19
0 327 317 316 315 337 336 335 334 277
0
0 0 4704 0
4 QDFF
-14 -44 14 -36
3 U95
-11 -46 10 -38
0
15 DVCC=16;DGND=8;
85 %D [%16bi %8bi %1i %2i %3i %4i %9i]
+ [%16bo %1o %2o %3o %4o %9o %5o %6o %7o %8o] %M
0
11 typeDigital
5 DIP16
19

0 1 2 3 4 5 6 7 8 9
1 2 3 4 5 6 7 8 9 0
65 0 0 0 1 0 0 0
1 U
5368 0 0
2
5.89979e-315 5.50703e-315
0
5 4011~
219 2511 2138 0 3 22
0 329 328 294
0
0 0 608 0
4 4011
-7 -24 21 -16
5 U118A
-18 -12 17 -4
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 9 0
65 0 0 0 4 1 42 0
1 U
8293 0 0
2
5.89979e-315 5.50833e-315
0
5 4011~
219 2516 1989 0 3 22
0 330 329 296
0
0 0 608 0
4 4011
-7 -24 21 -16
4 U92D
-17 -9 11 -1
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 9 0
65 0 0 0 4 4 33 0
1 U
3232 0 0
2
5.89979e-315 5.50963e-315
0
5 4011~
219 2519 1810 0 3 22
0 328 330 303
0
0 0 608 0
4 4011
-7 -24 21 -16
4 U92C
-21 -13 7 -5
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 8 9 10 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 9 0
65 0 0 0 4 3 33 0
1 U
6644 0 0
2
5.89979e-315 5.51092e-315
0
4 4008
219 2272 2216 0 14 29
0 13 14 15 16 221 220 219 218 642
281 280 279 278 300
0
0 0 4832 0
4 4008
-14 -60 14 -52
4 U113
-14 -61 14 -53
0
15 DVDD=16;DGND=8;
126 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 1 3 5 7 15 2 4 6 9
10 11 12 13 14 1 3 5 7 15
2 4 6 9 10 11 12 13 14 0
65 0 0 512 1 0 0 0
1 U
4978 0 0
2
5.89979e-315 5.51222e-315
0
14 Logic Display~
6 2360 2169 0 1 2
10 300
0
0 0 53872 512
6 100MEG
3 -16 45 -8
4 L133
-14 -21 14 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
9207 0 0
2
5.89979e-315 5.51286e-315
0
14 Logic Display~
6 2436 2170 0 1 2
10 281
0
0 0 53872 512
6 100MEG
3 -16 45 -8
4 L134
-14 -21 14 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
6998 0 0
2
5.89979e-315 5.51351e-315
0
14 Logic Display~
6 2423 2170 0 1 2
10 280
0
0 0 53872 512
6 100MEG
3 -16 45 -8
4 L135
-14 -21 14 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3175 0 0
2
5.89979e-315 5.51416e-315
0
14 Logic Display~
6 2410 2169 0 1 2
10 279
0
0 0 53872 512
6 100MEG
3 -16 45 -8
4 L136
-14 -21 14 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3378 0 0
2
5.89979e-315 5.51481e-315
0
14 Logic Display~
6 2397 2169 0 1 2
10 278
0
0 0 53872 512
6 100MEG
3 -16 45 -8
4 L137
-14 -21 14 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
922 0 0
2
5.89979e-315 5.51545e-315
0
4 4008
219 2272 2050 0 14 29
0 225 224 223 222 221 220 219 218 643
285 284 283 282 301
0
0 0 4832 0
4 4008
-14 -60 14 -52
4 U116
-14 -61 14 -53
0
15 DVDD=16;DGND=8;
126 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 1 3 5 7 15 2 4 6 9
10 11 12 13 14 1 3 5 7 15
2 4 6 9 10 11 12 13 14 0
65 0 0 512 1 0 0 0
1 U
6891 0 0
2
5.89979e-315 5.5161e-315
0
14 Logic Display~
6 2360 2003 0 1 2
10 301
0
0 0 53872 512
6 100MEG
3 -16 45 -8
4 L138
-14 -21 14 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
5407 0 0
2
5.89979e-315 5.51675e-315
0
14 Logic Display~
6 2436 2003 0 1 2
10 285
0
0 0 53872 512
6 100MEG
3 -16 45 -8
4 L139
-14 -21 14 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
7349 0 0
2
5.89979e-315 5.5174e-315
0
14 Logic Display~
6 2423 2004 0 1 2
10 284
0
0 0 53872 512
6 100MEG
3 -16 45 -8
4 L140
-14 -21 14 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3919 0 0
2
5.89979e-315 5.51804e-315
0
14 Logic Display~
6 2410 2004 0 1 2
10 283
0
0 0 53872 512
6 100MEG
3 -16 45 -8
4 L141
-14 -21 14 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
9747 0 0
2
5.89979e-315 5.51869e-315
0
14 Logic Display~
6 2397 2004 0 1 2
10 282
0
0 0 53872 512
6 100MEG
3 -16 45 -8
4 L142
-14 -21 14 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
5310 0 0
2
5.89979e-315 5.51934e-315
0
14 Logic Display~
6 2396 1846 0 1 2
10 311
0
0 0 53872 512
6 100MEG
3 -16 45 -8
4 L147
-14 -21 14 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
4318 0 0
2
5.89979e-315 5.51999e-315
0
14 Logic Display~
6 2409 1846 0 1 2
10 312
0
0 0 53872 512
6 100MEG
3 -16 45 -8
4 L146
-14 -21 14 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3917 0 0
2
5.89979e-315 5.52063e-315
0
14 Logic Display~
6 2422 1846 0 1 2
10 313
0
0 0 53872 512
6 100MEG
3 -16 45 -8
4 L145
-14 -21 14 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
7930 0 0
2
5.89979e-315 5.52128e-315
0
14 Logic Display~
6 2435 1846 0 1 2
10 314
0
0 0 53872 512
6 100MEG
3 -16 45 -8
4 L144
-14 -21 14 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
6128 0 0
2
5.89979e-315 5.52193e-315
0
14 Logic Display~
6 2359 1844 0 1 2
10 302
0
0 0 53872 512
6 100MEG
3 -16 45 -8
4 L143
-14 -21 14 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
7346 0 0
2
5.89979e-315 5.52258e-315
0
4 4008
219 2271 1889 0 14 29
0 13 14 15 16 225 224 223 222 644
314 313 312 311 302
0
0 0 4832 0
4 4008
-14 -60 14 -52
4 U114
-14 -61 14 -53
0
15 DVDD=16;DGND=8;
126 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 1 3 5 7 15 2 4 6 9
10 11 12 13 14 1 3 5 7 15
2 4 6 9 10 11 12 13 14 0
65 0 0 512 1 0 0 0
1 U
8577 0 0
2
5.89979e-315 5.52322e-315
0
9 Inverter~
13 1126 1555 0 2 22
0 343 344
0
0 0 608 180
6 74LS04
-21 -19 21 -11
5 U110D
-12 -20 23 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 9 8 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 4 39 0
1 U
3372 0 0
2
5.89979e-315 5.52387e-315
0
8 2-In OR~
219 861 1604 0 3 22
0 344 346 391
0
0 0 608 0
6 74LS32
-21 -24 21 -16
5 U111A
-11 -14 24 -6
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 40 0
1 U
3741 0 0
2
5.89979e-315 5.52452e-315
0
8 2-In OR~
219 863 1566 0 3 22
0 345 344 392
0
0 0 608 0
6 74LS32
-21 -24 21 -16
5 U100D
-8 -13 27 -5
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 38 0
1 U
5813 0 0
2
5.89979e-315 5.52517e-315
0
14 Logic Display~
6 1841 2012 0 1 2
10 351
0
0 0 53872 512
6 100MEG
3 -16 45 -8
4 L121
-14 -21 14 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3213 0 0
2
5.89979e-315 5.52581e-315
0
14 Logic Display~
6 1828 2012 0 1 2
10 350
0
0 0 53872 512
6 100MEG
3 -16 45 -8
4 L122
-14 -21 14 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3694 0 0
2
5.89979e-315 5.52646e-315
0
14 Logic Display~
6 1815 2012 0 1 2
10 349
0
0 0 53872 512
6 100MEG
3 -16 45 -8
4 L123
-14 -21 14 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
4327 0 0
2
5.89979e-315 5.52711e-315
0
14 Logic Display~
6 1802 2012 0 1 2
10 348
0
0 0 53872 512
6 100MEG
3 -16 45 -8
4 L124
-14 -21 14 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
8800 0 0
2
5.89979e-315 5.52776e-315
0
14 Logic Display~
6 1465 2011 0 1 2
10 352
0
0 0 53872 512
6 100MEG
3 -16 45 -8
4 L132
-14 -21 14 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3406 0 0
2
5.89979e-315 5.52841e-315
0
14 Logic Display~
6 1478 2011 0 1 2
10 353
0
0 0 53872 512
6 100MEG
3 -16 45 -8
4 L131
-14 -21 14 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
6455 0 0
2
5.89979e-315 5.52905e-315
0
14 Logic Display~
6 1491 2011 0 1 2
10 354
0
0 0 53872 512
6 100MEG
3 -16 45 -8
4 L130
-14 -21 14 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
9319 0 0
2
5.89979e-315 5.5297e-315
0
14 Logic Display~
6 1504 2011 0 1 2
10 355
0
0 0 53872 512
6 100MEG
3 -16 45 -8
4 L129
-14 -21 14 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3172 0 0
2
5.89979e-315 5.53035e-315
0
14 Logic Display~
6 1157 2010 0 1 2
10 359
0
0 0 53872 512
6 100MEG
3 -16 45 -8
4 L120
-14 -21 14 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
38 0 0
2
5.89979e-315 5.531e-315
0
14 Logic Display~
6 1144 2010 0 1 2
10 358
0
0 0 53872 512
6 100MEG
3 -16 45 -8
4 L119
-14 -21 14 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
376 0 0
2
5.89979e-315 5.53164e-315
0
14 Logic Display~
6 1131 2010 0 1 2
10 357
0
0 0 53872 512
6 100MEG
3 -16 45 -8
4 L118
-14 -21 14 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
6666 0 0
2
5.89979e-315 5.53229e-315
0
14 Logic Display~
6 1118 2010 0 1 2
10 356
0
0 0 53872 512
6 100MEG
3 -16 45 -8
4 L117
-14 -21 14 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
9365 0 0
2
5.89979e-315 5.53294e-315
0
9 Inverter~
13 1547 1841 0 2 22
0 364 361
0
0 0 608 270
6 74LS04
-21 -19 21 -11
5 U110C
-15 -15 20 -7
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 5 6 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 3 39 0
1 U
3251 0 0
2
5.89979e-315 5.53359e-315
0
9 Inverter~
13 1260 1826 0 2 22
0 366 362
0
0 0 608 270
6 74LS04
-21 -19 21 -11
5 U110B
-8 -5 27 3
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 3 4 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 2 39 0
1 U
5481 0 0
2
5.89979e-315 5.53423e-315
0
9 Inverter~
13 898 1809 0 2 22
0 365 363
0
0 0 608 270
6 74LS04
-21 -19 21 -11
5 U110A
-13 -12 22 -4
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 1 39 0
1 U
7788 0 0
2
5.89979e-315 5.53488e-315
0
9 8-In NOR~
219 1858 2245 0 9 19
0 341 339 338 260 255 201 198 645 367
0
0 0 608 90
4 4078
-7 -24 21 -16
4 U109
-5 -15 23 -7
0
15 DVDD=14;DGND=7;
97 %D [%14bi %7bi %1i %2i %3i %4i %5i %6i %7i %8i]
+ [%14bo %1o %2o %3o %4o %5o %6o %7o %8o %9o] %M
0
12 type:digital
5 DIP14
19

0 2 3 4 5 9 10 11 12 13
2 3 4 5 9 10 11 12 13 0
65 0 0 512 1 0 0 0
1 U
3273 0 0
2
5.89979e-315 5.53553e-315
0
9 8-In NOR~
219 1509 2240 0 9 19
0 347 340 339 275 260 226 201 199 368
0
0 0 608 90
4 4078
-7 -24 21 -16
4 U108
-11 -17 17 -9
0
15 DVDD=14;DGND=7;
97 %D [%14bi %7bi %1i %2i %3i %4i %5i %6i %7i %8i]
+ [%14bo %1o %2o %3o %4o %5o %6o %7o %8o %9o] %M
0
12 type:digital
5 DIP14
19

0 2 3 4 5 9 10 11 12 13
2 3 4 5 9 10 11 12 13 0
65 0 0 0 1 0 0 0
1 U
3761 0 0
2
5.89979e-315 5.53618e-315
0
9 8-In NOR~
219 1168 2236 0 9 19
0 360 340 338 275 255 226 200 17 369
0
0 0 608 90
4 4078
-7 -24 21 -16
4 U101
-6 -15 22 -7
0
15 DVDD=14;DGND=7;
97 %D [%14bi %7bi %1i %2i %3i %4i %5i %6i %7i %8i]
+ [%14bo %1o %2o %3o %4o %5o %6o %7o %8o %9o] %M
0
12 type:digital
5 DIP14
19

0 2 3 4 5 9 10 11 12 13
2 3 4 5 9 10 11 12 13 0
65 0 0 0 1 0 0 0
1 U
3226 0 0
2
5.89979e-315 5.53682e-315
0
9 Inverter~
13 1053 2253 0 2 22
0 373 372
0
0 0 608 90
6 74LS04
-21 -19 21 -11
4 U91D
-12 3 16 11
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 9 8 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 4 32 0
1 U
4244 0 0
2
44286.3 201
0
9 8-In NOR~
219 1050 2309 0 9 19
0 363 341 77 646 647 648 649 650 373
0
0 0 608 90
4 4078
-7 -24 21 -16
4 U106
-8 -16 20 -8
0
15 DVDD=14;DGND=7;
97 %D [%14bi %7bi %1i %2i %3i %4i %5i %6i %7i %8i]
+ [%14bo %1o %2o %3o %4o %5o %6o %7o %8o %9o] %M
0
12 type:digital
5 DIP14
19

0 2 3 4 5 9 10 11 12 13
2 3 4 5 9 10 11 12 13 0
65 0 0 512 1 0 0 0
1 U
5225 0 0
2
44286.3 202
0
9 Inverter~
13 1744 2264 0 2 22
0 374 370
0
0 0 608 90
6 74LS04
-21 -19 21 -11
4 U91F
-7 0 21 8
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 13 12 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 6 32 0
1 U
768 0 0
2
44286.3 203
0
9 8-In NOR~
219 1741 2320 0 9 19
0 361 347 651 652 653 654 655 656 374
0
0 0 608 90
4 4078
-7 -24 21 -16
4 U107
-4 -17 24 -9
0
15 DVDD=14;DGND=7;
97 %D [%14bi %7bi %1i %2i %3i %4i %5i %6i %7i %8i]
+ [%14bo %1o %2o %3o %4o %5o %6o %7o %8o %9o] %M
0
12 type:digital
5 DIP14
19

0 2 3 4 5 9 10 11 12 13
2 3 4 5 9 10 11 12 13 0
65 0 0 512 1 0 0 0
1 U
5735 0 0
2
44286.3 204
0
9 Inverter~
13 1402 2254 0 2 22
0 375 371
0
0 0 608 90
6 74LS04
-21 -19 21 -11
4 U91E
-9 0 19 8
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 11 10 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 5 32 0
1 U
5881 0 0
2
44286.3 205
0
9 8-In NOR~
219 1399 2310 0 9 19
0 362 360 657 658 659 660 661 662 375
0
0 0 608 90
4 4078
-7 -24 21 -16
4 U105
-8 -14 20 -6
0
15 DVDD=14;DGND=7;
97 %D [%14bi %7bi %1i %2i %3i %4i %5i %6i %7i %8i]
+ [%14bo %1o %2o %3o %4o %5o %6o %7o %8o %9o] %M
0
12 type:digital
5 DIP14
19

0 2 3 4 5 9 10 11 12 13
2 3 4 5 9 10 11 12 13 0
65 0 0 512 1 0 0 0
1 U
3275 0 0
2
44286.3 206
0
10 Buffer 3S~
219 1782 2164 0 3 22
0 342 370 376
0
0 0 608 602
8 BUFFER3S
-27 -51 29 -43
5 U104A
11 -5 46 3
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
0
22

0 2 1 3 2 1 3 5 4 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 26 0
1 U
4203 0 0
2
44286.3 207
0
10 Buffer 3S~
219 1447 2151 0 3 22
0 342 371 377
0
0 0 608 602
8 BUFFER3S
-27 -51 29 -43
4 U12A
-11 0 17 8
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
0
22

0 2 1 3 2 1 3 5 4 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 25 0
1 U
3440 0 0
2
44286.3 208
0
10 Buffer 3S~
219 1097 2161 0 3 22
0 342 372 378
0
0 0 608 602
8 BUFFER3S
-27 -51 29 -43
4 U82D
-15 2 13 10
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
0
22

0 12 13 11 2 1 3 5 4 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 27 0
1 U
9102 0 0
2
44286.3 209
0
13 Quad 3-State~
48 1864 2074 0 9 19
0 351 350 349 348 218 219 220 221 367
0
0 0 4704 0
8 QUAD3STA
-28 -44 28 -36
4 U103
-14 -46 14 -38
0
15 DVCC=16;DGND=8;
85 %D [%16bi %8bi %1i %2i %3i %4i %9i]
+ [%16bo %1o %2o %3o %4o %9o %5o %6o %7o %8o] %M
0
12 type:digital
5 DIP16
19

0 1 2 3 4 5 6 7 8 9
1 2 3 4 5 6 7 8 9 0
65 0 0 0 1 0 0 0
1 U
5586 0 0
2
44286.3 210
0
13 Quad 3-State~
48 1528 2076 0 9 19
0 355 354 353 352 222 223 224 225 368
0
0 0 4704 0
8 QUAD3STA
-28 -44 28 -36
3 U81
-11 -46 10 -38
0
15 DVCC=16;DGND=8;
85 %D [%16bi %8bi %1i %2i %3i %4i %9i]
+ [%16bo %1o %2o %3o %4o %9o %5o %6o %7o %8o] %M
0
12 type:digital
5 DIP16
19

0 1 2 3 4 5 6 7 8 9
1 2 3 4 5 6 7 8 9 0
65 0 0 0 1 0 0 0
1 U
525 0 0
2
44286.3 211
0
13 Quad 3-State~
48 1174 2079 0 9 19
0 359 358 357 356 16 15 14 13 369
0
0 0 4704 0
8 QUAD3STA
-28 -44 28 -36
4 U102
-14 -46 14 -38
0
15 DVCC=16;DGND=8;
85 %D [%16bi %8bi %1i %2i %3i %4i %9i]
+ [%16bo %1o %2o %3o %4o %9o %5o %6o %7o %8o] %M
0
12 type:digital
5 DIP16
19

0 1 2 3 4 5 6 7 8 9
1 2 3 4 5 6 7 8 9 0
65 0 0 0 1 0 0 0
1 U
6206 0 0
2
44286.3 212
0
14 Logic Display~
6 1542 1623 0 1 2
10 387
0
0 0 53872 602
6 100MEG
3 -16 45 -8
3 L22
13 -1 34 7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3418 0 0
2
5.89979e-315 5.53747e-315
0
14 Logic Display~
6 1455 1625 0 1 2
10 388
0
0 0 53872 602
6 100MEG
3 -16 45 -8
3 L21
13 -1 34 7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
9312 0 0
2
5.89979e-315 5.53812e-315
0
14 Logic Display~
6 1371 1622 0 1 2
10 389
0
0 0 53872 602
6 100MEG
3 -16 45 -8
3 L18
13 -1 34 7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
7419 0 0
2
5.89979e-315 5.53877e-315
0
14 Logic Display~
6 1274 1624 0 1 2
10 390
0
0 0 53872 602
6 100MEG
3 -16 45 -8
3 L17
13 -1 34 7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
472 0 0
2
5.89979e-315 5.53941e-315
0
9 Inverter~
13 964 1568 0 2 22
0 392 395
0
0 0 608 0
6 74LS04
-21 -19 21 -11
4 U74F
-7 -15 21 -7
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 13 12 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 6 19 0
1 U
4714 0 0
2
5.89979e-315 5.54006e-315
0
9 Inverter~
13 964 1586 0 2 22
0 391 394
0
0 0 608 0
6 74LS04
-21 -19 21 -11
4 U91A
-8 -11 20 -3
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 1 32 0
1 U
9386 0 0
2
5.89979e-315 5.54071e-315
0
9 Inverter~
13 966 1608 0 2 22
0 392 393
0
0 0 608 0
6 74LS04
-21 -19 21 -11
4 U91B
-4 -9 24 -1
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 3 4 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 2 32 0
1 U
7610 0 0
2
5.89979e-315 5.54136e-315
0
9 Inverter~
13 964 1668 0 2 22
0 391 396
0
0 0 608 0
6 74LS04
-21 -19 21 -11
4 U91C
-6 -14 22 -6
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 5 6 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 3 32 0
1 U
3482 0 0
2
5.89979e-315 5.542e-315
0
5 4011~
219 1014 1577 0 3 22
0 395 394 365
0
0 0 608 0
4 4011
-7 -24 21 -16
4 U89D
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 9 0
65 0 0 0 4 4 31 0
1 U
3608 0 0
2
5.89979e-315 5.54265e-315
0
5 4011~
219 1013 1617 0 3 22
0 393 391 366
0
0 0 608 0
4 4011
-7 -24 21 -16
4 U92A
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 9 0
65 0 0 0 4 1 33 0
1 U
6397 0 0
2
5.89979e-315 5.5433e-315
0
5 4011~
219 1014 1659 0 3 22
0 392 396 364
0
0 0 608 0
4 4011
-7 -24 21 -16
4 U92B
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 5 6 4 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 9 0
65 0 0 0 4 2 33 0
1 U
3967 0 0
2
5.89979e-315 5.54395e-315
0
12 Quad D Flop~
47 1097 2079 0 9 19
0 400 399 398 397 359 358 357 356 378
0
0 0 4704 0
4 QDFF
-14 -44 14 -36
3 U11
-11 -46 10 -38
0
15 DVCC=16;DGND=8;
85 %D [%16bi %8bi %1i %2i %3i %4i %9i]
+ [%16bo %1o %2o %3o %4o %9o %5o %6o %7o %8o] %M
0
11 typeDigital
5 DIP16
19

0 1 2 3 4 5 6 7 8 9
1 2 3 4 5 6 7 8 9 0
65 0 0 0 1 0 0 0
1 U
8621 0 0
2
5.89979e-315 5.54459e-315
0
12 Quad D Flop~
47 1447 2076 0 9 19
0 408 407 406 405 355 354 353 352 377
0
0 0 4704 0
4 QDFF
-14 -44 14 -36
3 U13
-11 -46 10 -38
0
15 DVCC=16;DGND=8;
85 %D [%16bi %8bi %1i %2i %3i %4i %9i]
+ [%16bo %1o %2o %3o %4o %9o %5o %6o %7o %8o] %M
0
11 typeDigital
5 DIP16
19

0 1 2 3 4 5 6 7 8 9
1 2 3 4 5 6 7 8 9 0
65 0 0 0 1 0 0 0
1 U
8901 0 0
2
5.89979e-315 5.54524e-315
0
12 Quad D Flop~
47 1781 2074 0 9 19
0 404 403 402 401 351 350 349 348 376
0
0 0 4704 0
4 QDFF
-14 -44 14 -36
3 U83
-11 -46 10 -38
0
15 DVCC=16;DGND=8;
85 %D [%16bi %8bi %1i %2i %3i %4i %9i]
+ [%16bo %1o %2o %3o %4o %9o %5o %6o %7o %8o] %M
0
11 typeDigital
5 DIP16
19

0 1 2 3 4 5 6 7 8 9
1 2 3 4 5 6 7 8 9 0
65 0 0 0 1 0 0 0
1 U
7385 0 0
2
5.89979e-315 5.54589e-315
0
8 2-In OR~
219 1333 2002 0 3 22
0 386 16 408
0
0 0 608 0
6 74LS32
-21 -24 21 -16
4 U84D
-4 -9 24 -1
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 28 0
1 U
6519 0 0
2
5.89979e-315 5.54654e-315
0
8 2-In OR~
219 1334 2049 0 3 22
0 385 15 407
0
0 0 608 0
6 74LS32
-21 -24 21 -16
4 U85A
-7 -12 21 -4
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 29 0
1 U
552 0 0
2
5.89979e-315 5.54719e-315
0
8 2-In OR~
219 1333 2096 0 3 22
0 384 14 406
0
0 0 608 0
6 74LS32
-21 -24 21 -16
4 U85B
-6 -9 22 -1
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 29 0
1 U
5551 0 0
2
5.89979e-315 5.54783e-315
0
8 2-In OR~
219 1333 2144 0 3 22
0 383 13 405
0
0 0 608 0
6 74LS32
-21 -24 21 -16
4 U85C
-6 -10 22 -2
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 9 10 8 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 29 0
1 U
8715 0 0
2
5.89979e-315 5.54848e-315
0
8 2-In OR~
219 1685 2004 0 3 22
0 382 222 404
0
0 0 608 0
6 74LS32
-21 -24 21 -16
4 U85D
-6 -9 22 -1
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 29 0
1 U
9763 0 0
2
5.89979e-315 5.54913e-315
0
8 2-In OR~
219 1684 2049 0 3 22
0 381 223 403
0
0 0 608 0
6 74LS32
-21 -24 21 -16
4 U86A
-8 -12 20 -4
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 30 0
1 U
8443 0 0
2
5.89979e-315 5.54978e-315
0
8 2-In OR~
219 1683 2088 0 3 22
0 380 224 402
0
0 0 608 0
6 74LS32
-21 -24 21 -16
4 U86B
-7 -13 21 -5
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 30 0
1 U
3719 0 0
2
5.89979e-315 5.55042e-315
0
8 2-In OR~
219 1682 2128 0 3 22
0 379 225 401
0
0 0 608 0
6 74LS32
-21 -24 21 -16
4 U86C
-7 -9 21 -1
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 9 10 8 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 30 0
1 U
8671 0 0
2
5.89979e-315 5.55107e-315
0
10 Buffer 3S~
219 1261 1603 0 3 22
0 412 343 390
0
0 0 608 270
8 BUFFER3S
-27 -51 29 -43
4 U79B
14 -5 42 3
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
0
22

0 5 4 6 2 1 3 5 4 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 23 0
1 U
7168 0 0
2
5.89979e-315 5.55172e-315
0
10 Buffer 3S~
219 1358 1600 0 3 22
0 411 343 389
0
0 0 608 270
8 BUFFER3S
-27 -51 29 -43
4 U80B
14 -5 42 3
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
0
22

0 5 4 6 2 1 3 5 4 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 24 0
1 U
49 0 0
2
5.89979e-315 5.55237e-315
0
10 Buffer 3S~
219 1441 1599 0 3 22
0 410 343 388
0
0 0 608 270
8 BUFFER3S
-27 -51 29 -43
4 U80C
14 -5 42 3
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
0
22

0 9 10 8 2 1 3 5 4 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 24 0
1 U
6536 0 0
2
5.89979e-315 5.55301e-315
0
10 Buffer 3S~
219 1529 1606 0 3 22
0 409 343 387
0
0 0 608 270
8 BUFFER3S
-27 -51 29 -43
4 U80D
14 -5 42 3
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
0
22

0 12 13 11 2 1 3 5 4 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 24 0
1 U
3931 0 0
2
5.89979e-315 5.55366e-315
0
13 Quad 3-State~
48 1604 1808 0 9 19
0 387 388 389 390 382 381 380 379 364
0
0 0 4704 270
8 QUAD3STA
-28 -44 28 -36
3 U88
42 -1 63 7
0
15 DVCC=16;DGND=8;
85 %D [%16bi %8bi %1i %2i %3i %4i %9i]
+ [%16bo %1o %2o %3o %4o %9o %5o %6o %7o %8o] %M
0
12 type:digital
5 DIP16
19

0 1 2 3 4 5 6 7 8 9
1 2 3 4 5 6 7 8 9 0
65 0 0 0 1 0 0 0
1 U
4390 0 0
2
5.89979e-315 5.55398e-315
0
13 Quad 3-State~
48 1338 1807 0 9 19
0 387 388 389 390 386 385 384 383 366
0
0 0 4704 270
8 QUAD3STA
-28 -44 28 -36
3 U87
42 -1 63 7
0
15 DVCC=16;DGND=8;
85 %D [%16bi %8bi %1i %2i %3i %4i %9i]
+ [%16bo %1o %2o %3o %4o %9o %5o %6o %7o %8o] %M
0
12 type:digital
5 DIP16
19

0 1 2 3 4 5 6 7 8 9
1 2 3 4 5 6 7 8 9 0
65 0 0 0 1 0 0 0
1 U
3242 0 0
2
5.89979e-315 5.55431e-315
0
13 Quad 3-State~
48 1065 1805 0 9 19
0 387 388 389 390 197 196 195 194 365
0
0 0 4704 270
8 QUAD3STA
-28 -44 28 -36
3 U90
42 -1 63 7
0
15 DVCC=16;DGND=8;
85 %D [%16bi %8bi %1i %2i %3i %4i %9i]
+ [%16bo %1o %2o %3o %4o %9o %5o %6o %7o %8o] %M
0
12 type:digital
5 DIP16
19

0 1 2 3 4 5 6 7 8 9
1 2 3 4 5 6 7 8 9 0
65 0 0 0 1 0 0 0
1 U
6760 0 0
2
5.89979e-315 5.55463e-315
0
7 Pulser~
4 638 2199 0 10 12
0 663 664 342 665 0 0 5 5 6
7
0
0 0 4640 0
0
2 V9
-7 -28 7 -20
0
0
0
0
0
4 SIP2
9

0 1 2 3 4 1 2 3 4 0
0 0 0 512 1 0 0 0
1 V
5760 0 0
2
44286.3 213
0
10 Buffer 3S~
219 823 1007 0 3 22
0 414 92 125
0
0 0 608 270
8 BUFFER3S
-27 -51 29 -43
4 U76C
-1 -4 27 4
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
0
22

0 9 10 8 2 1 3 5 4 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 20 0
1 U
3781 0 0
2
5.89979e-315 5.55496e-315
0
10 Buffer 3S~
219 860 1007 0 3 22
0 413 92 126
0
0 0 608 270
8 BUFFER3S
-27 -51 29 -43
4 U76B
-1 -4 27 4
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
0
22

0 5 4 6 2 1 3 5 4 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 20 0
1 U
8545 0 0
2
5.89979e-315 5.55528e-315
0
10 Buffer 3S~
219 784 1007 0 3 22
0 415 92 124
0
0 0 608 270
8 BUFFER3S
-27 -51 29 -43
4 U76A
-1 -4 27 4
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
0
22

0 2 1 3 2 1 3 5 4 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 20 0
1 U
9739 0 0
2
5.89979e-315 5.5556e-315
0
10 Buffer 3S~
219 747 1007 0 3 22
0 416 92 123
0
0 0 608 270
8 BUFFER3S
-27 -51 29 -43
4 U62D
-1 -4 27 4
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
0
22

0 12 13 11 2 1 3 5 4 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 16 0
1 U
388 0 0
2
5.89979e-315 5.55593e-315
0
14 Logic Display~
6 602 1649 0 1 2
10 198
0
0 0 53872 602
6 100MEG
3 -16 45 -8
4 L112
10 -1 38 7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
4595 0 0
2
5.89979e-315 5.55625e-315
0
14 Logic Display~
6 602 1633 0 1 2
10 102
0
0 0 53872 602
6 100MEG
3 -16 45 -8
4 L111
10 -1 38 7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3173 0 0
2
5.89979e-315 5.55657e-315
0
14 Logic Display~
6 601 1601 0 1 2
10 71
0
0 0 53872 602
6 100MEG
3 -16 45 -8
4 L110
10 -1 38 7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
9261 0 0
2
5.89979e-315 5.5569e-315
0
14 Logic Display~
6 602 1617 0 1 2
10 78
0
0 0 53872 602
6 100MEG
3 -16 45 -8
4 L109
10 -1 38 7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3494 0 0
2
5.89979e-315 5.55722e-315
0
14 Logic Display~
6 602 1714 0 1 2
10 255
0
0 0 53872 602
6 100MEG
3 -16 45 -8
4 L108
10 -1 38 7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
9101 0 0
2
5.89979e-315 5.55755e-315
0
14 Logic Display~
6 602 1698 0 1 2
10 226
0
0 0 53872 602
6 100MEG
3 -16 45 -8
4 L107
10 -1 38 7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
358 0 0
2
5.89979e-315 5.55787e-315
0
14 Logic Display~
6 601 1666 0 1 2
10 200
0
0 0 53872 602
6 100MEG
3 -16 45 -8
4 L106
10 -1 38 7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3726 0 0
2
5.89979e-315 5.55819e-315
0
14 Logic Display~
6 602 1682 0 1 2
10 201
0
0 0 53872 602
6 100MEG
3 -16 45 -8
4 L105
10 -1 38 7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
999 0 0
2
5.89979e-315 5.55852e-315
0
14 Logic Display~
6 602 1745 0 1 2
10 275
0
0 0 53872 602
6 100MEG
3 -16 45 -8
4 L104
9 -1 37 7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
8787 0 0
2
5.89979e-315 5.55884e-315
0
14 Logic Display~
6 602 1730 0 1 2
10 260
0
0 0 53872 602
6 100MEG
3 -16 45 -8
4 L103
9 -1 37 7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3348 0 0
2
5.89979e-315 5.55917e-315
0
14 Logic Display~
6 602 1761 0 1 2
10 338
0
0 0 53872 602
6 100MEG
3 -16 45 -8
3 L57
13 -1 34 7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3395 0 0
2
5.89979e-315 5.55949e-315
0
14 Logic Display~
6 602 1777 0 1 2
10 339
0
0 0 53872 602
6 100MEG
3 -16 45 -8
3 L56
13 -1 34 7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
7740 0 0
2
5.89979e-315 5.55981e-315
0
14 Logic Display~
6 602 1795 0 1 2
10 340
0
0 0 53872 602
6 100MEG
3 -16 45 -8
3 L24
13 -1 34 7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
6480 0 0
2
5.89979e-315 5.56014e-315
0
14 Logic Display~
6 602 1842 0 1 2
10 360
0
0 0 53872 602
6 100MEG
3 -16 45 -8
3 L23
13 -2 34 6
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
342 0 0
2
5.89979e-315 5.56046e-315
0
4 4514
219 417 1760 0 22 45
0 420 419 418 417 421 52 360 347 341
340 339 338 275 260 255 226 201 200 198
102 78 71
0
0 0 4832 0
4 4514
-14 -87 14 -79
3 U75
-11 -88 10 -80
0
16 DVDD=24;DGND=12;
155 %D [%24bi %12bi %1i %2i %3i %4i %5i %6i]
+ [%24bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o %15o %16o %17o %18o %19o %20o %21o %22o] %M
0
12 type:digital
5 DIP24
45

0 22 21 3 2 1 23 11 9 10
8 7 6 5 4 18 17 20 19 14
13 16 15 22 21 3 2 1 23 11
9 10 8 7 6 5 4 18 17 20
19 14 13 16 15 0
65 0 0 0 1 0 0 0
1 U
9953 0 0
2
5.89979e-315 5.56078e-315
0
14 Logic Display~
6 602 1825 0 1 2
10 347
0
0 0 53872 602
6 100MEG
3 -16 45 -8
3 L20
12 -1 33 7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
361 0 0
2
5.89979e-315 5.56111e-315
0
14 Logic Display~
6 602 1811 0 1 2
10 341
0
0 0 53872 602
6 100MEG
3 -16 45 -8
3 L19
12 0 33 8
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3343 0 0
2
5.89979e-315 5.56143e-315
0
14 Logic Display~
6 480 1421 0 1 2
10 420
0
0 0 53872 512
6 100MEG
3 -16 45 -8
3 H24
-11 -21 10 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
7923 0 0
2
5.89979e-315 5.56176e-315
0
14 Logic Display~
6 499 1421 0 1 2
10 419
0
0 0 53872 512
6 100MEG
3 -16 45 -8
3 H23
-11 -21 10 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
6174 0 0
2
5.89979e-315 5.56208e-315
0
14 Logic Display~
6 518 1421 0 1 2
10 418
0
0 0 53872 512
6 100MEG
3 -16 45 -8
3 H22
-11 -21 10 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
6692 0 0
2
5.89979e-315 5.5624e-315
0
14 Logic Display~
6 538 1421 0 1 2
10 417
0
0 0 53872 512
6 100MEG
3 -16 45 -8
3 H21
-11 -21 10 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
8790 0 0
2
5.89979e-315 5.56273e-315
0
14 Logic Display~
6 2922 1696 0 1 2
10 67
0
0 0 53872 512
6 100MEG
3 -16 45 -8
3 H19
-11 -21 10 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
4595 0 0
2
5.89979e-315 5.56305e-315
0
14 Logic Display~
6 2902 1696 0 1 2
10 68
0
0 0 53872 512
6 100MEG
3 -16 45 -8
2 H3
-8 -21 6 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
667 0 0
2
5.89979e-315 5.56337e-315
0
14 Logic Display~
6 2883 1696 0 1 2
10 69
0
0 0 53872 512
6 100MEG
3 -16 45 -8
2 H1
-8 -21 6 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
8743 0 0
2
5.89979e-315 5.5637e-315
0
12 Quad D Flop~
47 3080 1729 0 9 19
0 425 424 423 422 67 68 69 70 154
0
0 0 4704 180
4 QDFF
-14 -44 14 -36
3 U40
-11 40 10 48
0
15 DVCC=16;DGND=8;
85 %D [%16bi %8bi %1i %2i %3i %4i %9i]
+ [%16bo %1o %2o %3o %4o %9o %5o %6o %7o %8o] %M
0
11 typeDigital
5 DIP16
19

0 1 2 3 4 5 6 7 8 9
1 2 3 4 5 6 7 8 9 0
65 0 0 0 1 0 0 0
1 U
8298 0 0
2
5.89979e-315 5.56402e-315
0
14 Logic Display~
6 2864 1696 0 1 2
10 70
0
0 0 53872 512
6 100MEG
3 -16 45 -8
3 H20
-11 -21 10 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
313 0 0
2
5.89979e-315 5.56435e-315
0
9 Inverter~
13 3264 1484 0 2 22
0 428 429
0
0 0 608 0
6 74LS04
-21 -19 21 -11
4 U74A
-14 -20 14 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 1 19 0
1 U
7548 0 0
2
5.89979e-315 5.56467e-315
0
8 2-In OR~
219 3307 1625 0 3 22
0 429 430 425
0
0 0 608 270
6 74LS32
-21 -24 21 -16
4 U69B
-14 8 14 16
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 18 0
1 U
8973 0 0
2
5.89979e-315 5.56499e-315
0
9 Inverter~
13 3274 1578 0 2 22
0 426 430
0
0 0 608 0
6 74LS04
-21 -19 21 -11
4 U64F
-14 -20 14 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 13 12 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 6 17 0
1 U
9712 0 0
2
5.89979e-315 5.56532e-315
0
9 8-In NOR~
219 3213 1484 0 9 19
0 446 445 444 443 442 441 440 439 428
0
0 0 608 0
4 4078
-7 -24 21 -16
3 U73
1 4 22 12
0
15 DVDD=14;DGND=7;
97 %D [%14bi %7bi %1i %2i %3i %4i %5i %6i %7i %8i]
+ [%14bo %1o %2o %3o %4o %5o %6o %7o %8o %9o] %M
0
12 type:digital
5 DIP14
19

0 2 3 4 5 9 10 11 12 13
2 3 4 5 9 10 11 12 13 0
65 0 0 0 1 0 0 0
1 U
4518 0 0
2
5.89979e-315 5.56564e-315
0
9 8-In NOR~
219 3225 1578 0 9 19
0 438 437 436 435 434 433 432 431 426
0
0 0 608 0
4 4078
-7 -24 21 -16
3 U72
-2 1 19 9
0
15 DVDD=14;DGND=7;
97 %D [%14bi %7bi %1i %2i %3i %4i %5i %6i %7i %8i]
+ [%14bo %1o %2o %3o %4o %5o %6o %7o %8o %9o] %M
0
12 type:digital
5 DIP14
19

0 2 3 4 5 9 10 11 12 13
2 3 4 5 9 10 11 12 13 0
65 0 0 0 1 0 0 0
1 U
5596 0 0
2
5.89979e-315 5.56596e-315
0
9 8-In NOR~
219 3208 1336 0 9 19
0 457 456 435 455 454 453 452 451 427
0
0 0 608 0
4 4078
-7 -24 21 -16
3 U71
-2 1 19 9
0
15 DVDD=14;DGND=7;
97 %D [%14bi %7bi %1i %2i %3i %4i %5i %6i %7i %8i]
+ [%14bo %1o %2o %3o %4o %5o %6o %7o %8o %9o] %M
0
12 type:digital
5 DIP14
19

0 2 3 4 5 9 10 11 12 13
2 3 4 5 9 10 11 12 13 0
65 0 0 0 1 0 0 0
1 U
692 0 0
2
5.89979e-315 5.56629e-315
0
9 8-In NOR~
219 3193 1251 0 9 19
0 465 464 463 462 461 460 459 458 450
0
0 0 608 0
4 4078
-7 -24 21 -16
3 U70
1 4 22 12
0
15 DVDD=14;DGND=7;
97 %D [%14bi %7bi %1i %2i %3i %4i %5i %6i %7i %8i]
+ [%14bo %1o %2o %3o %4o %5o %6o %7o %8o %9o] %M
0
12 type:digital
5 DIP14
19

0 2 3 4 5 9 10 11 12 13
2 3 4 5 9 10 11 12 13 0
65 0 0 0 1 0 0 0
1 U
6258 0 0
2
5.89979e-315 5.56661e-315
0
9 Inverter~
13 3260 1336 0 2 22
0 427 449
0
0 0 608 0
6 74LS04
-21 -19 21 -11
4 U64E
-14 -20 14 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 11 10 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 5 17 0
1 U
5578 0 0
2
5.89979e-315 5.56694e-315
0
8 2-In OR~
219 3309 1363 0 3 22
0 448 449 424
0
0 0 608 270
6 74LS32
-21 -24 21 -16
4 U69A
-12 9 16 17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 18 0
1 U
8709 0 0
2
5.89979e-315 5.56726e-315
0
9 Inverter~
13 3245 1251 0 2 22
0 450 448
0
0 0 608 0
6 74LS04
-21 -19 21 -11
4 U64D
-14 -20 14 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 9 8 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 4 17 0
1 U
9131 0 0
2
5.89979e-315 5.56758e-315
0
9 Inverter~
13 3240 1037 0 2 22
0 469 466
0
0 0 608 0
6 74LS04
-21 -19 21 -11
4 U64C
-14 -20 14 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 5 6 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 3 17 0
1 U
3645 0 0
2
5.89979e-315 5.56791e-315
0
8 2-In OR~
219 3269 1139 0 3 22
0 466 467 423
0
0 0 608 270
6 74LS32
-21 -24 21 -16
3 U7D
-9 9 12 17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 6 0
1 U
7613 0 0
2
5.89979e-315 5.56823e-315
0
9 Inverter~
13 3239 1111 0 2 22
0 468 467
0
0 0 608 0
6 74LS04
-21 -19 21 -11
4 U64B
-14 -20 14 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 3 4 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 2 17 0
1 U
9467 0 0
2
5.89979e-315 5.56856e-315
0
9 8-In NOR~
219 3186 1037 0 9 19
0 470 471 472 473 474 475 476 477 469
0
0 0 608 0
4 4078
-7 -24 21 -16
3 U68
-2 0 19 8
0
15 DVDD=14;DGND=7;
97 %D [%14bi %7bi %1i %2i %3i %4i %5i %6i %7i %8i]
+ [%14bo %1o %2o %3o %4o %5o %6o %7o %8o %9o] %M
0
12 type:digital
5 DIP14
19

0 2 3 4 5 9 10 11 12 13
2 3 4 5 9 10 11 12 13 0
65 0 0 0 1 0 0 0
1 U
3932 0 0
2
5.89979e-315 5.56888e-315
0
9 8-In NOR~
219 3186 1111 0 9 19
0 478 479 480 447 481 482 483 484 468
0
0 0 608 0
4 4078
-7 -24 21 -16
3 U67
-2 1 19 9
0
15 DVDD=14;DGND=7;
97 %D [%14bi %7bi %1i %2i %3i %4i %5i %6i %7i %8i]
+ [%14bo %1o %2o %3o %4o %5o %6o %7o %8o %9o] %M
0
12 type:digital
5 DIP14
19

0 2 3 4 5 9 10 11 12 13
2 3 4 5 9 10 11 12 13 0
65 0 0 0 1 0 0 0
1 U
5288 0 0
2
5.89979e-315 5.5692e-315
0
9 8-In NOR~
219 3177 883 0 9 19
0 492 491 490 489 488 487 486 485 501
0
0 0 608 0
4 4078
-7 -24 21 -16
3 U66
-2 1 19 9
0
15 DVDD=14;DGND=7;
97 %D [%14bi %7bi %1i %2i %3i %4i %5i %6i %7i %8i]
+ [%14bo %1o %2o %3o %4o %5o %6o %7o %8o %9o] %M
0
12 type:digital
5 DIP14
19

0 2 3 4 5 9 10 11 12 13
2 3 4 5 9 10 11 12 13 0
65 0 0 0 1 0 0 0
1 U
4934 0 0
2
5.89979e-315 5.56953e-315
0
9 8-In NOR~
219 3177 811 0 9 19
0 500 499 498 497 496 495 494 493 503
0
0 0 608 0
4 4078
-7 -24 21 -16
3 U65
-2 0 19 8
0
15 DVDD=14;DGND=7;
97 %D [%14bi %7bi %1i %2i %3i %4i %5i %6i %7i %8i]
+ [%14bo %1o %2o %3o %4o %5o %6o %7o %8o %9o] %M
0
12 type:digital
5 DIP14
19

0 2 3 4 5 9 10 11 12 13
2 3 4 5 9 10 11 12 13 0
65 0 0 0 1 0 0 0
1 U
5987 0 0
2
5.89979e-315 5.56985e-315
0
9 Inverter~
13 3231 883 0 2 22
0 501 502
0
0 0 608 0
6 74LS04
-21 -19 21 -11
4 U64A
-14 -20 14 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 1 17 0
1 U
7737 0 0
2
5.89979e-315 5.57017e-315
0
8 2-In OR~
219 3258 907 0 3 22
0 504 502 422
0
0 0 608 270
6 74LS32
-21 -24 21 -16
3 U7C
-8 12 13 20
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 9 10 8 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 6 0
1 U
4200 0 0
2
5.89979e-315 5.5705e-315
0
9 Inverter~
13 3236 811 0 2 22
0 503 504
0
0 0 608 0
6 74LS04
-21 -19 21 -11
4 U56F
-14 -20 14 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 13 12 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 6 12 0
1 U
5780 0 0
2
5.89979e-315 5.57082e-315
0
7 Pulser~
4 1791 1670 0 10 12
0 666 667 153 668 0 0 5 5 6
7
0
0 0 4640 0
0
3 V26
-10 -28 11 -20
0
0
0
0
0
4 SIP2
9

0 1 2 3 4 1 2 3 4 0
0 0 0 512 1 0 0 0
1 V
6490 0 0
2
5.89979e-315 5.57115e-315
0
10 Buffer 3S~
219 3036 1215 0 3 22
0 153 166 505
0
0 0 608 512
8 BUFFER3S
-27 -51 29 -43
4 U62B
-14 -20 14 -12
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
0
22

0 5 4 6 2 1 3 5 4 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 16 0
1 U
8663 0 0
2
5.89979e-315 5.57147e-315
0
10 Buffer 3S~
219 2711 1216 0 3 22
0 153 168 506
0
0 0 608 512
8 BUFFER3S
-27 -51 29 -43
4 U62A
-14 -20 14 -12
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
0
22

0 2 1 3 2 1 3 5 4 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 16 0
1 U
318 0 0
2
5.89979e-315 5.57179e-315
0
10 Buffer 3S~
219 2424 1213 0 3 22
0 153 170 507
0
0 0 608 512
8 BUFFER3S
-27 -51 29 -43
4 U61D
-14 -20 14 -12
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
0
22

0 12 13 11 2 1 3 5 4 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 15 0
1 U
348 0 0
2
5.89979e-315 5.57212e-315
0
10 Buffer 3S~
219 2132 1215 0 3 22
0 153 172 508
0
0 0 608 512
8 BUFFER3S
-27 -51 29 -43
4 U61C
-14 -20 14 -12
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
0
22

0 9 10 8 2 1 3 5 4 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 15 0
1 U
8551 0 0
2
5.89979e-315 5.57244e-315
0
10 Buffer 3S~
219 3031 1447 0 3 22
0 153 158 509
0
0 0 608 512
8 BUFFER3S
-27 -51 29 -43
4 U61B
-14 -20 14 -12
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
0
22

0 5 4 6 2 1 3 5 4 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 15 0
1 U
7295 0 0
2
5.89979e-315 5.57276e-315
0
10 Buffer 3S~
219 2706 1449 0 3 22
0 153 160 510
0
0 0 608 512
8 BUFFER3S
-27 -51 29 -43
4 U61A
-14 -20 14 -12
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
0
22

0 2 1 3 2 1 3 5 4 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 15 0
1 U
9900 0 0
2
5.89979e-315 5.57309e-315
0
10 Buffer 3S~
219 2415 1449 0 3 22
0 153 162 511
0
0 0 608 512
8 BUFFER3S
-27 -51 29 -43
4 U60D
-14 -20 14 -12
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
0
22

0 12 13 11 2 1 3 5 4 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 14 0
1 U
8725 0 0
2
5.89979e-315 5.57341e-315
0
10 Buffer 3S~
219 2122 1450 0 3 22
0 153 164 512
0
0 0 608 512
8 BUFFER3S
-27 -51 29 -43
4 U60C
-14 -20 14 -12
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
0
22

0 9 10 8 2 1 3 5 4 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 14 0
1 U
366 0 0
2
5.89979e-315 5.57374e-315
0
10 Buffer 3S~
219 3038 999 0 3 22
0 153 174 513
0
0 0 608 512
8 BUFFER3S
-27 -51 29 -43
4 U60B
-14 -20 14 -12
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
0
22

0 5 4 6 2 1 3 5 4 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 14 0
1 U
5762 0 0
2
5.89979e-315 5.57406e-315
0
10 Buffer 3S~
219 2710 999 0 3 22
0 153 176 514
0
0 0 608 512
8 BUFFER3S
-27 -51 29 -43
4 U60A
-14 -20 14 -12
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
0
22

0 2 1 3 2 1 3 5 4 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 14 0
1 U
4943 0 0
2
5.89979e-315 5.57438e-315
0
10 Buffer 3S~
219 2426 996 0 3 22
0 153 178 515
0
0 0 608 512
8 BUFFER3S
-27 -51 29 -43
4 U59D
-14 -20 14 -12
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
0
22

0 12 13 11 2 1 3 5 4 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 13 0
1 U
3435 0 0
2
5.89979e-315 5.57471e-315
0
10 Buffer 3S~
219 2136 999 0 3 22
0 153 180 516
0
0 0 608 512
8 BUFFER3S
-27 -51 29 -43
4 U59C
-14 -20 14 -12
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
0
22

0 9 10 8 2 1 3 5 4 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 13 0
1 U
8705 0 0
2
5.89979e-315 5.57503e-315
0
10 Buffer 3S~
219 3025 777 0 3 22
0 153 182 517
0
0 0 608 512
8 BUFFER3S
-27 -51 29 -43
4 U59B
-14 -20 14 -12
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
0
22

0 5 4 6 2 1 3 5 4 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 13 0
1 U
4331 0 0
2
5.89979e-315 5.57535e-315
0
10 Buffer 3S~
219 2716 779 0 3 22
0 153 184 518
0
0 0 608 512
8 BUFFER3S
-27 -51 29 -43
4 U59A
-14 -20 14 -12
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
0
22

0 2 1 3 2 1 3 5 4 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 13 0
1 U
787 0 0
2
5.89979e-315 5.57568e-315
0
10 Buffer 3S~
219 2435 778 0 3 22
0 153 187 519
0
0 0 608 512
8 BUFFER3S
-27 -51 29 -43
4 U14D
-14 -20 14 -12
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
0
22

0 12 13 11 2 1 3 5 4 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 10 0
1 U
3655 0 0
2
5.89979e-315 5.576e-315
0
14 Logic Display~
6 2872 1462 0 1 2
10 525
0
0 0 53872 512
6 100MEG
3 -16 45 -8
3 H18
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
6682 0 0
2
5.89979e-315 5.57633e-315
0
14 Logic Display~
6 2887 1462 0 1 2
10 524
0
0 0 53872 512
6 100MEG
3 -16 45 -8
4 L102
-14 -21 14 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
582 0 0
2
5.89979e-315 5.57665e-315
0
14 Logic Display~
6 2901 1462 0 1 2
10 523
0
0 0 53872 512
6 100MEG
3 -16 45 -8
4 L101
-14 -21 14 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3125 0 0
2
5.89979e-315 5.57697e-315
0
14 Logic Display~
6 2915 1462 0 1 2
10 522
0
0 0 53872 512
6 100MEG
3 -16 45 -8
4 L100
-14 -21 14 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
5466 0 0
2
5.89979e-315 5.5773e-315
0
13 Quad 3-State~
48 2978 1518 0 9 19
0 525 524 523 522 485 484 451 431 521
0
0 0 4704 782
8 QUAD3STA
-28 -44 28 -36
3 U58
-64 -1 -43 7
0
15 DVCC=16;DGND=8;
85 %D [%16bi %8bi %1i %2i %3i %4i %9i]
+ [%16bo %1o %2o %3o %4o %9o %5o %6o %7o %8o] %M
0
12 type:digital
5 DIP16
19

0 1 2 3 4 5 6 7 8 9
1 2 3 4 5 6 7 8 9 0
65 0 0 0 1 0 0 0
1 U
52 0 0
2
5.89979e-315 5.57762e-315
0
9 Inverter~
13 3029 1521 0 2 22
0 157 521
0
0 0 608 180
6 74LS04
-21 -19 21 -11
4 U56B
-8 -20 20 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 3 4 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 2 12 0
1 U
3898 0 0
2
5.89979e-315 5.57795e-315
0
14 Logic Display~
6 2546 1464 0 1 2
10 530
0
0 0 53872 512
6 100MEG
3 -16 45 -8
3 H17
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
9413 0 0
2
5.89979e-315 5.57827e-315
0
14 Logic Display~
6 2561 1464 0 1 2
10 529
0
0 0 53872 512
6 100MEG
3 -16 45 -8
3 L99
-11 -21 10 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
8576 0 0
2
5.89979e-315 5.57859e-315
0
14 Logic Display~
6 2575 1464 0 1 2
10 528
0
0 0 53872 512
6 100MEG
3 -16 45 -8
3 L98
-11 -21 10 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
622 0 0
2
5.89979e-315 5.57892e-315
0
14 Logic Display~
6 2589 1464 0 1 2
10 527
0
0 0 53872 512
6 100MEG
3 -16 45 -8
3 L97
-11 -21 10 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
9152 0 0
2
5.89979e-315 5.57924e-315
0
13 Quad 3-State~
48 2652 1522 0 9 19
0 530 529 528 527 486 483 452 432 526
0
0 0 4704 782
8 QUAD3STA
-28 -44 28 -36
3 U57
-64 -1 -43 7
0
15 DVCC=16;DGND=8;
85 %D [%16bi %8bi %1i %2i %3i %4i %9i]
+ [%16bo %1o %2o %3o %4o %9o %5o %6o %7o %8o] %M
0
12 type:digital
5 DIP16
19

0 1 2 3 4 5 6 7 8 9
1 2 3 4 5 6 7 8 9 0
65 0 0 0 1 0 0 0
1 U
783 0 0
2
5.89979e-315 5.57956e-315
0
9 Inverter~
13 2703 1525 0 2 22
0 159 526
0
0 0 608 180
6 74LS04
-21 -19 21 -11
4 U56A
-8 -20 20 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 1 12 0
1 U
4262 0 0
2
5.89979e-315 5.57989e-315
0
14 Logic Display~
6 2258 1464 0 1 2
10 535
0
0 0 53872 512
6 100MEG
3 -16 45 -8
3 H16
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
6121 0 0
2
5.89979e-315 5.58021e-315
0
14 Logic Display~
6 2273 1464 0 1 2
10 534
0
0 0 53872 512
6 100MEG
3 -16 45 -8
3 L96
-11 -21 10 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3879 0 0
2
5.89979e-315 5.58054e-315
0
14 Logic Display~
6 2287 1464 0 1 2
10 533
0
0 0 53872 512
6 100MEG
3 -16 45 -8
3 L95
-11 -21 10 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
7345 0 0
2
5.89979e-315 5.58086e-315
0
14 Logic Display~
6 2301 1464 0 1 2
10 532
0
0 0 53872 512
6 100MEG
3 -16 45 -8
3 L94
-11 -21 10 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3198 0 0
2
5.89979e-315 5.58118e-315
0
13 Quad 3-State~
48 2364 1520 0 9 19
0 535 534 533 532 487 482 453 433 531
0
0 0 4704 782
8 QUAD3STA
-28 -44 28 -36
3 U55
-64 -1 -43 7
0
15 DVCC=16;DGND=8;
85 %D [%16bi %8bi %1i %2i %3i %4i %9i]
+ [%16bo %1o %2o %3o %4o %9o %5o %6o %7o %8o] %M
0
12 type:digital
5 DIP16
19

0 1 2 3 4 5 6 7 8 9
1 2 3 4 5 6 7 8 9 0
65 0 0 0 1 0 0 0
1 U
9849 0 0
2
5.89979e-315 5.58151e-315
0
9 Inverter~
13 2415 1523 0 2 22
0 161 531
0
0 0 608 180
6 74LS04
-21 -19 21 -11
4 U49F
-8 -20 20 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 13 12 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 6 11 0
1 U
479 0 0
2
5.89979e-315 5.58183e-315
0
14 Logic Display~
6 1967 1465 0 1 2
10 540
0
0 0 53872 512
6 100MEG
3 -16 45 -8
3 H15
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3905 0 0
2
5.89979e-315 5.58215e-315
0
14 Logic Display~
6 1982 1465 0 1 2
10 539
0
0 0 53872 512
6 100MEG
3 -16 45 -8
3 L93
-11 -21 10 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
4394 0 0
2
5.89979e-315 5.58248e-315
0
14 Logic Display~
6 1996 1465 0 1 2
10 538
0
0 0 53872 512
6 100MEG
3 -16 45 -8
3 L92
-11 -21 10 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
4391 0 0
2
5.89979e-315 5.5828e-315
0
14 Logic Display~
6 2010 1465 0 1 2
10 537
0
0 0 53872 512
6 100MEG
3 -16 45 -8
3 L91
-11 -21 10 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3681 0 0
2
5.89979e-315 5.58313e-315
0
13 Quad 3-State~
48 2073 1523 0 9 19
0 540 539 538 537 488 481 454 434 536
0
0 0 4704 782
8 QUAD3STA
-28 -44 28 -36
3 U54
-64 -1 -43 7
0
15 DVCC=16;DGND=8;
85 %D [%16bi %8bi %1i %2i %3i %4i %9i]
+ [%16bo %1o %2o %3o %4o %9o %5o %6o %7o %8o] %M
0
12 type:digital
5 DIP16
19

0 1 2 3 4 5 6 7 8 9
1 2 3 4 5 6 7 8 9 0
65 0 0 0 1 0 0 0
1 U
6466 0 0
2
5.89979e-315 5.58345e-315
0
9 Inverter~
13 2124 1526 0 2 22
0 163 536
0
0 0 608 180
6 74LS04
-21 -19 21 -11
4 U49E
-8 -20 20 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 11 10 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 5 11 0
1 U
5230 0 0
2
5.89979e-315 5.58377e-315
0
14 Logic Display~
6 2878 1230 0 1 2
10 545
0
0 0 53872 512
6 100MEG
3 -16 45 -8
3 H14
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
8324 0 0
2
5.89979e-315 5.5841e-315
0
14 Logic Display~
6 2893 1230 0 1 2
10 544
0
0 0 53872 512
6 100MEG
3 -16 45 -8
3 L90
-11 -21 10 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3445 0 0
2
5.89979e-315 5.58442e-315
0
14 Logic Display~
6 2907 1230 0 1 2
10 543
0
0 0 53872 512
6 100MEG
3 -16 45 -8
3 L89
-11 -21 10 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
7543 0 0
2
5.89979e-315 5.58474e-315
0
14 Logic Display~
6 2921 1230 0 1 2
10 542
0
0 0 53872 512
6 100MEG
3 -16 45 -8
3 L88
-11 -21 10 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
6187 0 0
2
5.89979e-315 5.58507e-315
0
13 Quad 3-State~
48 2984 1285 0 9 19
0 545 544 543 542 489 447 455 435 541
0
0 0 4704 782
8 QUAD3STA
-28 -44 28 -36
3 U53
-64 -1 -43 7
0
15 DVCC=16;DGND=8;
85 %D [%16bi %8bi %1i %2i %3i %4i %9i]
+ [%16bo %1o %2o %3o %4o %9o %5o %6o %7o %8o] %M
0
12 type:digital
5 DIP16
19

0 1 2 3 4 5 6 7 8 9
1 2 3 4 5 6 7 8 9 0
65 0 0 0 1 0 0 0
1 U
5476 0 0
2
5.89979e-315 5.58539e-315
0
9 Inverter~
13 3035 1288 0 2 22
0 165 541
0
0 0 608 180
6 74LS04
-21 -19 21 -11
4 U49D
-8 -20 20 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 9 8 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 4 11 0
1 U
3936 0 0
2
5.89979e-315 5.58572e-315
0
14 Logic Display~
6 2552 1231 0 1 2
10 550
0
0 0 53872 512
6 100MEG
3 -16 45 -8
3 H13
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
5770 0 0
2
5.89979e-315 5.58604e-315
0
14 Logic Display~
6 2567 1231 0 1 2
10 549
0
0 0 53872 512
6 100MEG
3 -16 45 -8
3 L87
-11 -21 10 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
7884 0 0
2
5.89979e-315 5.58636e-315
0
14 Logic Display~
6 2581 1231 0 1 2
10 548
0
0 0 53872 512
6 100MEG
3 -16 45 -8
3 L86
-11 -21 10 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3690 0 0
2
5.89979e-315 5.58669e-315
0
14 Logic Display~
6 2595 1231 0 1 2
10 547
0
0 0 53872 512
6 100MEG
3 -16 45 -8
3 L85
-11 -21 10 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3611 0 0
2
5.89979e-315 5.58701e-315
0
13 Quad 3-State~
48 2658 1287 0 9 19
0 550 549 548 547 490 480 435 436 546
0
0 0 4704 782
8 QUAD3STA
-28 -44 28 -36
3 U52
-64 -1 -43 7
0
15 DVCC=16;DGND=8;
85 %D [%16bi %8bi %1i %2i %3i %4i %9i]
+ [%16bo %1o %2o %3o %4o %9o %5o %6o %7o %8o] %M
0
12 type:digital
5 DIP16
19

0 1 2 3 4 5 6 7 8 9
1 2 3 4 5 6 7 8 9 0
65 0 0 0 1 0 0 0
1 U
7912 0 0
2
5.89979e-315 5.58734e-315
0
9 Inverter~
13 2709 1290 0 2 22
0 167 546
0
0 0 608 180
6 74LS04
-21 -19 21 -11
4 U49C
-8 -20 20 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 5 6 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 3 11 0
1 U
6416 0 0
2
5.89979e-315 5.58766e-315
0
14 Logic Display~
6 2264 1228 0 1 2
10 555
0
0 0 53872 512
6 100MEG
3 -16 45 -8
3 H12
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
7278 0 0
2
5.89979e-315 5.58798e-315
0
14 Logic Display~
6 2279 1228 0 1 2
10 554
0
0 0 53872 512
6 100MEG
3 -16 45 -8
3 L84
-11 -21 10 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
6804 0 0
2
5.89979e-315 5.58831e-315
0
14 Logic Display~
6 2293 1228 0 1 2
10 553
0
0 0 53872 512
6 100MEG
3 -16 45 -8
3 L83
-11 -21 10 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
9568 0 0
2
5.89979e-315 5.58863e-315
0
14 Logic Display~
6 2307 1228 0 1 2
10 552
0
0 0 53872 512
6 100MEG
3 -16 45 -8
3 L82
-11 -21 10 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
7178 0 0
2
5.89979e-315 5.58895e-315
0
13 Quad 3-State~
48 2370 1284 0 9 19
0 555 554 553 552 491 479 456 437 551
0
0 0 4704 782
8 QUAD3STA
-28 -44 28 -36
3 U51
-64 -1 -43 7
0
15 DVCC=16;DGND=8;
85 %D [%16bi %8bi %1i %2i %3i %4i %9i]
+ [%16bo %1o %2o %3o %4o %9o %5o %6o %7o %8o] %M
0
12 type:digital
5 DIP16
19

0 1 2 3 4 5 6 7 8 9
1 2 3 4 5 6 7 8 9 0
65 0 0 0 1 0 0 0
1 U
7982 0 0
2
5.89979e-315 5.58928e-315
0
9 Inverter~
13 2421 1287 0 2 22
0 169 551
0
0 0 608 180
6 74LS04
-21 -19 21 -11
4 U49B
-8 -20 20 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 3 4 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 2 11 0
1 U
513 0 0
2
5.89979e-315 5.5896e-315
0
14 Logic Display~
6 1973 1230 0 1 2
10 560
0
0 0 53872 512
6 100MEG
3 -16 45 -8
3 H11
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
8190 0 0
2
5.89979e-315 5.58993e-315
0
14 Logic Display~
6 1988 1230 0 1 2
10 559
0
0 0 53872 512
6 100MEG
3 -16 45 -8
3 L81
-11 -21 10 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
5209 0 0
2
5.89979e-315 5.59025e-315
0
14 Logic Display~
6 2002 1230 0 1 2
10 558
0
0 0 53872 512
6 100MEG
3 -16 45 -8
3 L80
-11 -21 10 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
7239 0 0
2
5.89979e-315 5.59057e-315
0
14 Logic Display~
6 2016 1230 0 1 2
10 557
0
0 0 53872 512
6 100MEG
3 -16 45 -8
3 L79
-11 -21 10 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
9474 0 0
2
5.89979e-315 5.5909e-315
0
13 Quad 3-State~
48 2079 1287 0 9 19
0 560 559 558 557 492 478 457 438 556
0
0 0 4704 782
8 QUAD3STA
-28 -44 28 -36
3 U50
-64 -1 -43 7
0
15 DVCC=16;DGND=8;
85 %D [%16bi %8bi %1i %2i %3i %4i %9i]
+ [%16bo %1o %2o %3o %4o %9o %5o %6o %7o %8o] %M
0
12 type:digital
5 DIP16
19

0 1 2 3 4 5 6 7 8 9
1 2 3 4 5 6 7 8 9 0
65 0 0 0 1 0 0 0
1 U
3783 0 0
2
5.89979e-315 5.59122e-315
0
9 Inverter~
13 2130 1290 0 2 22
0 171 556
0
0 0 608 180
6 74LS04
-21 -19 21 -11
4 U49A
-8 -20 20 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 1 11 0
1 U
5422 0 0
2
5.89979e-315 5.59154e-315
0
14 Logic Display~
6 2881 1014 0 1 2
10 565
0
0 0 53872 512
6 100MEG
3 -16 45 -8
3 H10
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
8527 0 0
2
5.89979e-315 5.59187e-315
0
14 Logic Display~
6 2896 1014 0 1 2
10 564
0
0 0 53872 512
6 100MEG
3 -16 45 -8
3 L78
-11 -21 10 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
761 0 0
2
5.89979e-315 5.59219e-315
0
14 Logic Display~
6 2910 1014 0 1 2
10 563
0
0 0 53872 512
6 100MEG
3 -16 45 -8
3 L77
-11 -21 10 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
7323 0 0
2
5.89979e-315 5.59252e-315
0
14 Logic Display~
6 2924 1014 0 1 2
10 562
0
0 0 53872 512
6 100MEG
3 -16 45 -8
3 L76
-11 -21 10 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
8543 0 0
2
5.89979e-315 5.59284e-315
0
13 Quad 3-State~
48 2987 1069 0 9 19
0 565 564 563 562 493 477 458 439 561
0
0 0 4704 782
8 QUAD3STA
-28 -44 28 -36
3 U48
-64 -1 -43 7
0
15 DVCC=16;DGND=8;
85 %D [%16bi %8bi %1i %2i %3i %4i %9i]
+ [%16bo %1o %2o %3o %4o %9o %5o %6o %7o %8o] %M
0
12 type:digital
5 DIP16
19

0 1 2 3 4 5 6 7 8 9
1 2 3 4 5 6 7 8 9 0
65 0 0 0 1 0 0 0
1 U
4240 0 0
2
5.89979e-315 5.59316e-315
0
9 Inverter~
13 3038 1072 0 2 22
0 173 561
0
0 0 608 180
6 74LS04
-21 -19 21 -11
4 U41F
-8 -20 20 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 13 12 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 6 8 0
1 U
7857 0 0
2
5.89979e-315 5.59349e-315
0
14 Logic Display~
6 2555 1014 0 1 2
10 570
0
0 0 53872 512
6 100MEG
3 -16 45 -8
2 H9
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
7255 0 0
2
5.89979e-315 5.59381e-315
0
14 Logic Display~
6 2570 1014 0 1 2
10 569
0
0 0 53872 512
6 100MEG
3 -16 45 -8
3 L75
-11 -21 10 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
7736 0 0
2
5.89979e-315 5.59413e-315
0
14 Logic Display~
6 2584 1014 0 1 2
10 568
0
0 0 53872 512
6 100MEG
3 -16 45 -8
3 L74
-11 -21 10 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
5435 0 0
2
5.89979e-315 5.59446e-315
0
14 Logic Display~
6 2598 1014 0 1 2
10 567
0
0 0 53872 512
6 100MEG
3 -16 45 -8
3 L73
-11 -21 10 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3446 0 0
2
5.89979e-315 5.59478e-315
0
13 Quad 3-State~
48 2661 1072 0 9 19
0 570 569 568 567 494 476 459 440 566
0
0 0 4704 782
8 QUAD3STA
-28 -44 28 -36
3 U47
-64 -1 -43 7
0
15 DVCC=16;DGND=8;
85 %D [%16bi %8bi %1i %2i %3i %4i %9i]
+ [%16bo %1o %2o %3o %4o %9o %5o %6o %7o %8o] %M
0
12 type:digital
5 DIP16
19

0 1 2 3 4 5 6 7 8 9
1 2 3 4 5 6 7 8 9 0
65 0 0 0 1 0 0 0
1 U
3914 0 0
2
5.89979e-315 5.59511e-315
0
9 Inverter~
13 2712 1075 0 2 22
0 175 566
0
0 0 608 180
6 74LS04
-21 -19 21 -11
4 U41E
-8 -20 20 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 11 10 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 5 8 0
1 U
3948 0 0
2
5.89979e-315 5.59527e-315
0
14 Logic Display~
6 2267 1010 0 1 2
10 575
0
0 0 53872 512
6 100MEG
3 -16 45 -8
2 H8
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3901 0 0
2
5.89979e-315 5.59543e-315
0
14 Logic Display~
6 2282 1010 0 1 2
10 574
0
0 0 53872 512
6 100MEG
3 -16 45 -8
3 L72
-11 -21 10 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
6295 0 0
2
5.89979e-315 5.59559e-315
0
14 Logic Display~
6 2296 1010 0 1 2
10 573
0
0 0 53872 512
6 100MEG
3 -16 45 -8
3 L71
-11 -21 10 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
332 0 0
2
5.89979e-315 5.59575e-315
0
14 Logic Display~
6 2310 1010 0 1 2
10 572
0
0 0 53872 512
6 100MEG
3 -16 45 -8
3 L70
-11 -21 10 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
9737 0 0
2
5.89979e-315 5.59592e-315
0
13 Quad 3-State~
48 2373 1067 0 9 19
0 575 574 573 572 495 475 460 441 571
0
0 0 4704 782
8 QUAD3STA
-28 -44 28 -36
3 U46
-64 -1 -43 7
0
15 DVCC=16;DGND=8;
85 %D [%16bi %8bi %1i %2i %3i %4i %9i]
+ [%16bo %1o %2o %3o %4o %9o %5o %6o %7o %8o] %M
0
12 type:digital
5 DIP16
19

0 1 2 3 4 5 6 7 8 9
1 2 3 4 5 6 7 8 9 0
65 0 0 0 1 0 0 0
1 U
9910 0 0
2
5.89979e-315 5.59608e-315
0
9 Inverter~
13 2424 1070 0 2 22
0 177 571
0
0 0 608 180
6 74LS04
-21 -19 21 -11
4 U41D
-8 -20 20 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 9 8 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 4 8 0
1 U
3834 0 0
2
5.89979e-315 5.59624e-315
0
14 Logic Display~
6 1976 1014 0 1 2
10 580
0
0 0 53872 512
6 100MEG
3 -16 45 -8
2 H7
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3138 0 0
2
5.89979e-315 5.5964e-315
0
14 Logic Display~
6 1991 1014 0 1 2
10 579
0
0 0 53872 512
6 100MEG
3 -16 45 -8
3 L69
-11 -21 10 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
5409 0 0
2
5.89979e-315 5.59656e-315
0
14 Logic Display~
6 2005 1014 0 1 2
10 578
0
0 0 53872 512
6 100MEG
3 -16 45 -8
3 L68
-11 -21 10 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
983 0 0
2
5.89979e-315 5.59673e-315
0
14 Logic Display~
6 2019 1014 0 1 2
10 577
0
0 0 53872 512
6 100MEG
3 -16 45 -8
3 L67
-11 -21 10 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
6652 0 0
2
5.89979e-315 5.59689e-315
0
13 Quad 3-State~
48 2082 1072 0 9 19
0 580 579 578 577 496 474 461 442 576
0
0 0 4704 782
8 QUAD3STA
-28 -44 28 -36
3 U45
-64 -1 -43 7
0
15 DVCC=16;DGND=8;
85 %D [%16bi %8bi %1i %2i %3i %4i %9i]
+ [%16bo %1o %2o %3o %4o %9o %5o %6o %7o %8o] %M
0
12 type:digital
5 DIP16
19

0 1 2 3 4 5 6 7 8 9
1 2 3 4 5 6 7 8 9 0
65 0 0 0 1 0 0 0
1 U
4281 0 0
2
5.89979e-315 5.59705e-315
0
9 Inverter~
13 2133 1075 0 2 22
0 179 576
0
0 0 608 180
6 74LS04
-21 -19 21 -11
4 U41C
-8 -20 20 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 5 6 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 3 8 0
1 U
6847 0 0
2
5.89979e-315 5.59721e-315
0
14 Logic Display~
6 2871 790 0 1 2
10 584
0
0 0 53872 512
6 100MEG
3 -16 45 -8
2 H6
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
6543 0 0
2
5.89979e-315 5.59737e-315
0
14 Logic Display~
6 2886 790 0 1 2
10 583
0
0 0 53872 512
6 100MEG
3 -16 45 -8
3 L66
-11 -21 10 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
7168 0 0
2
5.89979e-315 5.59753e-315
0
14 Logic Display~
6 2900 790 0 1 2
10 582
0
0 0 53872 512
6 100MEG
3 -16 45 -8
3 L65
-11 -21 10 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3828 0 0
2
5.89979e-315 5.5977e-315
0
14 Logic Display~
6 2914 790 0 1 2
10 581
0
0 0 53872 512
6 100MEG
3 -16 45 -8
3 L64
-11 -21 10 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
955 0 0
2
5.89979e-315 5.59786e-315
0
13 Quad 3-State~
48 2977 845 0 9 19
0 584 583 582 581 497 473 462 443 585
0
0 0 4704 782
8 QUAD3STA
-28 -44 28 -36
3 U43
-64 -1 -43 7
0
15 DVCC=16;DGND=8;
85 %D [%16bi %8bi %1i %2i %3i %4i %9i]
+ [%16bo %1o %2o %3o %4o %9o %5o %6o %7o %8o] %M
0
12 type:digital
5 DIP16
19

0 1 2 3 4 5 6 7 8 9
1 2 3 4 5 6 7 8 9 0
65 0 0 0 1 0 0 0
1 U
7782 0 0
2
5.89979e-315 5.59802e-315
0
9 Inverter~
13 3028 848 0 2 22
0 181 585
0
0 0 608 180
6 74LS04
-21 -19 21 -11
4 U41B
-8 -20 20 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 3 4 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 2 8 0
1 U
824 0 0
2
5.89979e-315 5.59818e-315
0
14 Logic Display~
6 2557 793 0 1 2
10 590
0
0 0 53872 512
6 100MEG
3 -16 45 -8
2 H5
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
6983 0 0
2
5.89979e-315 5.59834e-315
0
14 Logic Display~
6 2572 793 0 1 2
10 589
0
0 0 53872 512
6 100MEG
3 -16 45 -8
3 L63
-11 -21 10 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3185 0 0
2
5.89979e-315 5.59851e-315
0
14 Logic Display~
6 2586 793 0 1 2
10 588
0
0 0 53872 512
6 100MEG
3 -16 45 -8
3 L62
-11 -21 10 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
4213 0 0
2
5.89979e-315 5.59867e-315
0
14 Logic Display~
6 2600 793 0 1 2
10 587
0
0 0 53872 512
6 100MEG
3 -16 45 -8
3 L61
-11 -21 10 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
9765 0 0
2
5.89979e-315 5.59883e-315
0
13 Quad 3-State~
48 2663 851 0 9 19
0 590 589 588 587 498 472 463 444 586
0
0 0 4704 782
8 QUAD3STA
-28 -44 28 -36
3 U42
-64 -1 -43 7
0
15 DVCC=16;DGND=8;
85 %D [%16bi %8bi %1i %2i %3i %4i %9i]
+ [%16bo %1o %2o %3o %4o %9o %5o %6o %7o %8o] %M
0
12 type:digital
5 DIP16
19

0 1 2 3 4 5 6 7 8 9
1 2 3 4 5 6 7 8 9 0
65 0 0 0 1 0 0 0
1 U
8986 0 0
2
5.89979e-315 5.59899e-315
0
9 Inverter~
13 2714 854 0 2 22
0 183 586
0
0 0 608 180
6 74LS04
-21 -19 21 -11
4 U41A
-8 -20 20 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 1 8 0
1 U
3273 0 0
2
5.89979e-315 5.59915e-315
0
14 Logic Display~
6 2276 792 0 1 2
10 595
0
0 0 53872 512
6 100MEG
3 -16 45 -8
2 H2
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
5636 0 0
2
5.89979e-315 5.59932e-315
0
14 Logic Display~
6 2291 792 0 1 2
10 594
0
0 0 53872 512
6 100MEG
3 -16 45 -8
3 L54
-11 -21 10 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
327 0 0
2
5.89979e-315 5.59948e-315
0
14 Logic Display~
6 2305 792 0 1 2
10 593
0
0 0 53872 512
6 100MEG
3 -16 45 -8
3 L53
-11 -21 10 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
9233 0 0
2
5.89979e-315 5.59964e-315
0
14 Logic Display~
6 2319 792 0 1 2
10 592
0
0 0 53872 512
6 100MEG
3 -16 45 -8
3 L49
-11 -21 10 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3875 0 0
2
5.89979e-315 5.5998e-315
0
13 Quad 3-State~
48 2382 847 0 9 19
0 595 594 593 592 499 471 464 445 591
0
0 0 4704 782
8 QUAD3STA
-28 -44 28 -36
3 U39
-64 -1 -43 7
0
15 DVCC=16;DGND=8;
85 %D [%16bi %8bi %1i %2i %3i %4i %9i]
+ [%16bo %1o %2o %3o %4o %9o %5o %6o %7o %8o] %M
0
12 type:digital
5 DIP16
19

0 1 2 3 4 5 6 7 8 9
1 2 3 4 5 6 7 8 9 0
65 0 0 0 1 0 0 0
1 U
9991 0 0
2
5.89979e-315 5.59996e-315
0
9 Inverter~
13 2433 850 0 2 22
0 186 591
0
0 0 608 180
6 74LS04
-21 -19 21 -11
3 U2F
-5 -20 16 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 13 12 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 6 1 0
1 U
3221 0 0
2
5.89979e-315 5.60012e-315
0
14 Logic Display~
6 1975 796 0 1 2
10 599
0
0 0 53872 512
6 100MEG
3 -16 45 -8
2 H4
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
8874 0 0
2
5.89979e-315 5.60029e-315
0
14 Logic Display~
6 1990 796 0 1 2
10 598
0
0 0 53872 512
6 100MEG
3 -16 45 -8
3 L58
-11 -21 10 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
7400 0 0
2
5.89979e-315 5.60045e-315
0
14 Logic Display~
6 2004 796 0 1 2
10 597
0
0 0 53872 512
6 100MEG
3 -16 45 -8
3 L59
-11 -21 10 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3623 0 0
2
5.89979e-315 5.60061e-315
0
14 Logic Display~
6 2018 796 0 1 2
10 596
0
0 0 53872 512
6 100MEG
3 -16 45 -8
3 L60
-11 -21 10 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3311 0 0
2
5.89979e-315 5.60077e-315
0
13 Quad 3-State~
48 2081 853 0 9 19
0 599 598 597 596 500 470 465 446 600
0
0 0 4704 782
8 QUAD3STA
-28 -44 28 -36
3 U38
-64 -1 -43 7
0
15 DVCC=16;DGND=8;
85 %D [%16bi %8bi %1i %2i %3i %4i %9i]
+ [%16bo %1o %2o %3o %4o %9o %5o %6o %7o %8o] %M
0
12 type:digital
5 DIP16
19

0 1 2 3 4 5 6 7 8 9
1 2 3 4 5 6 7 8 9 0
65 0 0 0 1 0 0 0
1 U
5736 0 0
2
5.89979e-315 5.60093e-315
0
9 Inverter~
13 2132 856 0 2 22
0 185 600
0
0 0 608 180
6 74LS04
-21 -19 21 -11
3 U2E
-5 -20 16 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 11 10 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 5 1 0
1 U
3143 0 0
2
5.89979e-315 5.6011e-315
0
10 Buffer 3S~
219 2137 783 0 3 22
0 153 188 520
0
0 0 608 512
8 BUFFER3S
-27 -51 29 -43
4 U14C
-14 -20 14 -12
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
0
22

0 9 10 8 2 1 3 5 4 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 10 0
1 U
5835 0 0
2
5.89979e-315 5.60126e-315
0
13 Quad 3-State~
48 673 1086 0 9 19
0 611 610 609 608 126 125 124 123 92
0
0 0 4704 0
8 QUAD3STA
-28 -44 28 -36
3 U36
-11 -46 10 -38
0
15 DVCC=16;DGND=8;
85 %D [%16bi %8bi %1i %2i %3i %4i %9i]
+ [%16bo %1o %2o %3o %4o %9o %5o %6o %7o %8o] %M
0
12 type:digital
5 DIP16
19

0 1 2 3 4 5 6 7 8 9
1 2 3 4 5 6 7 8 9 0
65 0 0 0 1 0 0 0
1 U
5108 0 0
2
44286.3 214
0
12 Quad D Flop~
47 2984 999 0 9 19
0 604 603 602 601 565 564 563 562 513
0
0 0 4704 782
4 QDFF
-14 -44 14 -36
3 U34
-61 -4 -40 4
0
15 DVCC=16;DGND=8;
85 %D [%16bi %8bi %1i %2i %3i %4i %9i]
+ [%16bo %1o %2o %3o %4o %9o %5o %6o %7o %8o] %M
0
11 typeDigital
5 DIP16
19

0 1 2 3 4 5 6 7 8 9
1 2 3 4 5 6 7 8 9 0
65 0 0 0 1 0 0 0
1 U
3320 0 0
2
44286.3 215
0
12 Quad D Flop~
47 2981 1215 0 9 19
0 604 603 602 601 545 544 543 542 505
0
0 0 4704 782
4 QDFF
-14 -44 14 -36
3 U31
-61 -4 -40 4
0
15 DVCC=16;DGND=8;
85 %D [%16bi %8bi %1i %2i %3i %4i %9i]
+ [%16bo %1o %2o %3o %4o %9o %5o %6o %7o %8o] %M
0
11 typeDigital
5 DIP16
19

0 1 2 3 4 5 6 7 8 9
1 2 3 4 5 6 7 8 9 0
65 0 0 0 1 0 0 0
1 U
523 0 0
2
44286.3 216
0
12 Quad D Flop~
47 2975 1447 0 9 19
0 604 603 602 601 525 524 523 522 509
0
0 0 4704 782
4 QDFF
-14 -44 14 -36
3 U30
-61 -4 -40 4
0
15 DVCC=16;DGND=8;
85 %D [%16bi %8bi %1i %2i %3i %4i %9i]
+ [%16bo %1o %2o %3o %4o %9o %5o %6o %7o %8o] %M
0
11 typeDigital
5 DIP16
19

0 1 2 3 4 5 6 7 8 9
1 2 3 4 5 6 7 8 9 0
65 0 0 0 1 0 0 0
1 U
3557 0 0
2
44286.3 217
0
12 Quad D Flop~
47 2658 999 0 9 19
0 604 603 602 601 570 569 568 567 514
0
0 0 4704 782
4 QDFF
-14 -44 14 -36
3 U29
-61 -4 -40 4
0
15 DVCC=16;DGND=8;
85 %D [%16bi %8bi %1i %2i %3i %4i %9i]
+ [%16bo %1o %2o %3o %4o %9o %5o %6o %7o %8o] %M
0
11 typeDigital
5 DIP16
19

0 1 2 3 4 5 6 7 8 9
1 2 3 4 5 6 7 8 9 0
65 0 0 0 1 0 0 0
1 U
7246 0 0
2
44286.3 218
0
12 Quad D Flop~
47 2655 1216 0 9 19
0 604 603 602 601 550 549 548 547 506
0
0 0 4704 782
4 QDFF
-14 -44 14 -36
3 U27
-61 -4 -40 4
0
15 DVCC=16;DGND=8;
85 %D [%16bi %8bi %1i %2i %3i %4i %9i]
+ [%16bo %1o %2o %3o %4o %9o %5o %6o %7o %8o] %M
0
11 typeDigital
5 DIP16
19

0 1 2 3 4 5 6 7 8 9
1 2 3 4 5 6 7 8 9 0
65 0 0 0 1 0 0 0
1 U
3916 0 0
2
44286.3 219
0
12 Quad D Flop~
47 2649 1449 0 9 19
0 604 603 602 601 530 529 528 527 510
0
0 0 4704 782
4 QDFF
-14 -44 14 -36
3 U26
-61 -4 -40 4
0
15 DVCC=16;DGND=8;
85 %D [%16bi %8bi %1i %2i %3i %4i %9i]
+ [%16bo %1o %2o %3o %4o %9o %5o %6o %7o %8o] %M
0
11 typeDigital
5 DIP16
19

0 1 2 3 4 5 6 7 8 9
1 2 3 4 5 6 7 8 9 0
65 0 0 0 1 0 0 0
1 U
614 0 0
2
44286.3 220
0
12 Quad D Flop~
47 2370 996 0 9 19
0 604 603 602 601 575 574 573 572 515
0
0 0 4704 782
4 QDFF
-14 -44 14 -36
3 U25
-61 -4 -40 4
0
15 DVCC=16;DGND=8;
85 %D [%16bi %8bi %1i %2i %3i %4i %9i]
+ [%16bo %1o %2o %3o %4o %9o %5o %6o %7o %8o] %M
0
11 typeDigital
5 DIP16
19

0 1 2 3 4 5 6 7 8 9
1 2 3 4 5 6 7 8 9 0
65 0 0 0 1 0 0 0
1 U
8494 0 0
2
44286.3 221
0
12 Quad D Flop~
47 2367 1213 0 9 19
0 604 603 602 601 555 554 553 552 507
0
0 0 4704 782
4 QDFF
-14 -44 14 -36
3 U24
-61 -4 -40 4
0
15 DVCC=16;DGND=8;
85 %D [%16bi %8bi %1i %2i %3i %4i %9i]
+ [%16bo %1o %2o %3o %4o %9o %5o %6o %7o %8o] %M
0
11 typeDigital
5 DIP16
19

0 1 2 3 4 5 6 7 8 9
1 2 3 4 5 6 7 8 9 0
65 0 0 0 1 0 0 0
1 U
774 0 0
2
44286.3 222
0
12 Quad D Flop~
47 2361 1449 0 9 19
0 604 603 602 601 535 534 533 532 511
0
0 0 4704 782
4 QDFF
-14 -44 14 -36
3 U23
-61 -4 -40 4
0
15 DVCC=16;DGND=8;
85 %D [%16bi %8bi %1i %2i %3i %4i %9i]
+ [%16bo %1o %2o %3o %4o %9o %5o %6o %7o %8o] %M
0
11 typeDigital
5 DIP16
19

0 1 2 3 4 5 6 7 8 9
1 2 3 4 5 6 7 8 9 0
65 0 0 0 1 0 0 0
1 U
715 0 0
2
44286.3 223
0
12 Quad D Flop~
47 2070 1450 0 9 19
0 604 603 602 601 540 539 538 537 512
0
0 0 4704 782
4 QDFF
-14 -44 14 -36
3 U22
-61 -4 -40 4
0
15 DVCC=16;DGND=8;
85 %D [%16bi %8bi %1i %2i %3i %4i %9i]
+ [%16bo %1o %2o %3o %4o %9o %5o %6o %7o %8o] %M
0
11 typeDigital
5 DIP16
19

0 1 2 3 4 5 6 7 8 9
1 2 3 4 5 6 7 8 9 0
65 0 0 0 1 0 0 0
1 U
3281 0 0
2
44286.3 224
0
12 Quad D Flop~
47 2076 1215 0 9 19
0 604 603 602 601 560 559 558 557 508
0
0 0 4704 782
4 QDFF
-14 -44 14 -36
3 U21
-61 -4 -40 4
0
15 DVCC=16;DGND=8;
85 %D [%16bi %8bi %1i %2i %3i %4i %9i]
+ [%16bo %1o %2o %3o %4o %9o %5o %6o %7o %8o] %M
0
11 typeDigital
5 DIP16
19

0 1 2 3 4 5 6 7 8 9
1 2 3 4 5 6 7 8 9 0
65 0 0 0 1 0 0 0
1 U
3593 0 0
2
44286.3 225
0
12 Quad D Flop~
47 2079 999 0 9 19
0 604 603 602 601 580 579 578 577 516
0
0 0 4704 782
4 QDFF
-14 -44 14 -36
3 U18
-61 -4 -40 4
0
15 DVCC=16;DGND=8;
85 %D [%16bi %8bi %1i %2i %3i %4i %9i]
+ [%16bo %1o %2o %3o %4o %9o %5o %6o %7o %8o] %M
0
11 typeDigital
5 DIP16
19

0 1 2 3 4 5 6 7 8 9
1 2 3 4 5 6 7 8 9 0
65 0 0 0 1 0 0 0
1 U
7233 0 0
2
44286.3 226
0
12 Quad D Flop~
47 2974 777 0 9 19
0 604 603 602 601 584 583 582 581 517
0
0 0 4704 782
4 QDFF
-14 -44 14 -36
3 U17
-61 -4 -40 4
0
15 DVCC=16;DGND=8;
85 %D [%16bi %8bi %1i %2i %3i %4i %9i]
+ [%16bo %1o %2o %3o %4o %9o %5o %6o %7o %8o] %M
0
11 typeDigital
5 DIP16
19

0 1 2 3 4 5 6 7 8 9
1 2 3 4 5 6 7 8 9 0
65 0 0 0 1 0 0 0
1 U
3410 0 0
2
44286.3 227
0
12 Quad D Flop~
47 2660 779 0 9 19
0 604 603 602 601 590 589 588 587 518
0
0 0 4704 782
4 QDFF
-14 -44 14 -36
3 U16
-61 -4 -40 4
0
15 DVCC=16;DGND=8;
85 %D [%16bi %8bi %1i %2i %3i %4i %9i]
+ [%16bo %1o %2o %3o %4o %9o %5o %6o %7o %8o] %M
0
11 typeDigital
5 DIP16
19

0 1 2 3 4 5 6 7 8 9
1 2 3 4 5 6 7 8 9 0
65 0 0 0 1 0 0 0
1 U
3616 0 0
2
44286.3 228
0
12 Quad D Flop~
47 2379 778 0 9 19
0 604 603 602 601 595 594 593 592 519
0
0 0 4704 782
4 QDFF
-14 -44 14 -36
3 U15
-61 -4 -40 4
0
15 DVCC=16;DGND=8;
85 %D [%16bi %8bi %1i %2i %3i %4i %9i]
+ [%16bo %1o %2o %3o %4o %9o %5o %6o %7o %8o] %M
0
11 typeDigital
5 DIP16
19

0 1 2 3 4 5 6 7 8 9
1 2 3 4 5 6 7 8 9 0
65 0 0 0 1 0 0 0
1 U
5202 0 0
2
44286.3 229
0
10 Buffer 3S~
219 2202 579 0 3 22
0 605 90 603
0
0 0 608 0
8 BUFFER3S
-27 -51 29 -43
4 U14A
-14 -20 14 -12
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
0
22

0 2 1 3 2 1 3 5 4 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 10 0
1 U
9145 0 0
2
44286.3 230
0
14 Logic Display~
6 2217 1598 0 1 2
10 603
0
0 0 53872 692
6 100MEG
3 -16 45 -8
3 L42
11 0 32 8
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
9815 0 0
2
44286.3 231
0
10 Buffer 3S~
219 2495 584 0 3 22
0 606 90 602
0
0 0 608 0
8 BUFFER3S
-27 -51 29 -43
4 U32D
-14 -20 14 -12
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
0
22

0 12 13 11 2 1 3 5 4 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 9 0
1 U
4766 0 0
2
44286.3 232
0
14 Logic Display~
6 2510 1603 0 1 2
10 602
0
0 0 53872 692
6 100MEG
3 -16 45 -8
3 L45
11 0 32 8
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
8325 0 0
2
44286.3 233
0
10 Buffer 3S~
219 2798 590 0 3 22
0 91 90 601
0
0 0 608 0
8 BUFFER3S
-27 -51 29 -43
4 U32C
-14 -20 14 -12
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
0
22

0 9 10 8 2 1 3 5 4 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 9 0
1 U
7196 0 0
2
44286.3 234
0
14 Logic Display~
6 2813 1609 0 1 2
10 601
0
0 0 53872 692
6 100MEG
3 -16 45 -8
3 L44
11 0 32 8
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3567 0 0
2
44286.3 235
0
14 Logic Display~
6 1933 1604 0 1 2
10 604
0
0 0 53872 692
6 100MEG
3 -16 45 -8
3 L41
11 0 32 8
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
5877 0 0
2
44286.3 236
0
12 Quad D Flop~
47 2078 783 0 9 19
0 604 603 602 601 599 598 597 596 520
0
0 0 4704 782
4 QDFF
-14 -44 14 -36
3 U20
14 -26 35 -18
0
15 DVCC=16;DGND=8;
85 %D [%16bi %8bi %1i %2i %3i %4i %9i]
+ [%16bo %1o %2o %3o %4o %9o %5o %6o %7o %8o] %M
0
11 typeDigital
5 DIP16
19

0 1 2 3 4 5 6 7 8 9
1 2 3 4 5 6 7 8 9 0
65 0 0 0 1 0 0 0
1 U
4785 0 0
2
44286.3 237
0
10 Buffer 3S~
219 1917 584 0 3 22
0 607 90 604
0
0 0 608 0
8 BUFFER3S
-27 -51 29 -43
4 U32A
-14 -20 14 -12
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
0
22

0 2 1 3 2 1 3 5 4 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 9 0
1 U
3822 0 0
2
44286.3 238
0
12 Quad D Flop~
47 527 1086 0 9 19
0 76 75 74 73 611 610 609 608 132
0
0 0 4704 0
4 QDFF
-14 -44 14 -36
3 U19
-11 -46 10 -38
0
15 DVCC=16;DGND=8;
85 %D [%16bi %8bi %1i %2i %3i %4i %9i]
+ [%16bo %1o %2o %3o %4o %9o %5o %6o %7o %8o] %M
0
11 typeDigital
5 DIP16
19

0 1 2 3 4 5 6 7 8 9
1 2 3 4 5 6 7 8 9 0
65 0 0 0 1 0 0 0
1 U
7640 0 0
2
5.89979e-315 5.60142e-315
0
12 Quad D Flop~
47 579 1455 0 9 19
0 67 68 69 70 417 418 419 420 189
0
0 0 4704 180
4 QDFF
-14 -44 14 -36
3 U44
-11 40 10 48
0
15 DVCC=16;DGND=8;
85 %D [%16bi %8bi %1i %2i %3i %4i %9i]
+ [%16bo %1o %2o %3o %4o %9o %5o %6o %7o %8o] %M
0
11 typeDigital
5 DIP16
19

0 1 2 3 4 5 6 7 8 9
1 2 3 4 5 6 7 8 9 0
65 0 0 0 1 0 0 0
1 U
9221 0 0
2
5.89979e-315 5.60158e-315
0
7 Pulser~
4 315 1310 0 10 12
0 669 670 132 671 0 0 5 5 6
7
0
0 0 4640 0
0
2 V7
-7 -28 7 -20
0
0
0
0
0
4 SIP2
9

0 1 2 3 4 1 2 3 4 0
0 0 0 512 1 0 0 0
1 V
6484 0 0
2
44286.3 239
0
4 4514
219 1345 1088 0 30 45
0 119 120 121 122 155 156 185 186 183
181 179 177 175 173 171 169 167 165 163
161 159 157 0 0 0 0 0 0 0
3
0
0 0 4832 692
4 4514
-14 -87 14 -79
3 U33
-11 -88 10 -80
0
16 DVDD=24;DGND=12;
155 %D [%24bi %12bi %1i %2i %3i %4i %5i %6i]
+ [%24bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o %15o %16o %17o %18o %19o %20o %21o %22o] %M
0
12 type:digital
5 DIP24
45

0 22 21 3 2 1 23 11 9 10
8 7 6 5 4 18 17 20 19 14
13 16 15 22 21 3 2 1 23 11
9 10 8 7 6 5 4 18 17 20
19 14 13 16 15 0
65 0 0 0 1 0 0 0
1 U
3689 0 0
2
44286.3 240
0
14 Logic Display~
6 1465 1133 0 1 2
10 161
0
0 0 53872 602
6 100MEG
3 -16 45 -8
3 L25
12 0 33 8
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3952 0 0
2
44286.3 241
0
14 Logic Display~
6 1465 1147 0 1 2
10 159
0
0 0 53872 602
6 100MEG
3 -16 45 -8
3 L26
12 -1 33 7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3631 0 0
2
44286.3 242
0
14 Logic Display~
6 1465 1164 0 1 2
10 157
0
0 0 53872 602
6 100MEG
3 -16 45 -8
3 L27
13 -2 34 6
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
9359 0 0
2
44286.3 243
0
14 Logic Display~
6 1465 1117 0 1 2
10 163
0
0 0 53872 602
6 100MEG
3 -16 45 -8
3 L28
13 -1 34 7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
5584 0 0
2
44286.3 244
0
14 Logic Display~
6 1465 1099 0 1 2
10 165
0
0 0 53872 602
6 100MEG
3 -16 45 -8
3 L29
13 -1 34 7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
4973 0 0
2
44286.3 245
0
14 Logic Display~
6 1465 1083 0 1 2
10 167
0
0 0 53872 602
6 100MEG
3 -16 45 -8
3 L30
13 -1 34 7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3239 0 0
2
44286.3 246
0
14 Logic Display~
6 1465 1052 0 1 2
10 171
0
0 0 53872 602
6 100MEG
3 -16 45 -8
3 L31
13 -1 34 7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
4244 0 0
2
44286.3 247
0
14 Logic Display~
6 1465 1067 0 1 2
10 169
0
0 0 53872 602
6 100MEG
3 -16 45 -8
3 L32
13 -1 34 7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3391 0 0
2
44286.3 248
0
14 Logic Display~
6 1465 1004 0 1 2
10 177
0
0 0 53872 602
6 100MEG
3 -16 45 -8
3 L33
13 -1 34 7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
4243 0 0
2
44286.3 249
0
14 Logic Display~
6 1464 988 0 1 2
10 179
0
0 0 53872 602
6 100MEG
3 -16 45 -8
3 L34
13 -1 34 7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3907 0 0
2
44286.3 250
0
14 Logic Display~
6 1465 1020 0 1 2
10 175
0
0 0 53872 602
6 100MEG
3 -16 45 -8
3 L35
13 -1 34 7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
728 0 0
2
44286.3 251
0
14 Logic Display~
6 1465 1036 0 1 2
10 173
0
0 0 53872 602
6 100MEG
3 -16 45 -8
3 L36
14 -1 35 7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3585 0 0
2
44286.3 252
0
14 Logic Display~
6 1465 939 0 1 2
10 186
0
0 0 53872 602
6 100MEG
3 -16 45 -8
3 L37
13 -1 34 7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3565 0 0
2
44286.3 253
0
14 Logic Display~
6 1464 923 0 1 2
10 185
0
0 0 53872 602
6 100MEG
3 -16 45 -8
3 L38
13 -1 34 7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3966 0 0
2
44286.3 254
0
14 Logic Display~
6 1465 955 0 1 2
10 183
0
0 0 53872 602
6 100MEG
3 -16 45 -8
3 L39
13 -1 34 7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3714 0 0
2
44286.3 255
0
14 Logic Display~
6 1465 971 0 1 2
10 181
0
0 0 53872 602
6 100MEG
3 -16 45 -8
3 L40
13 -1 34 7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3406 0 0
2
44286.3 256
0
1203
3 1 2 0 0 12416 0 23 108 0 0 6
909 1395
924 1395
924 1430
1285 1430
1285 1311
1317 1311
2 0 3 0 0 4096 0 23 0 0 228 4
863 1404
820 1404
820 1433
815 1433
3 1 4 0 0 4224 0 93 23 0 0 4
809 1380
855 1380
855 1386
863 1386
1 5 5 0 0 8320 0 24 35 0 0 3
1288 782
1288 761
1316 761
2 5 6 0 0 4224 0 24 30 0 0 2
1279 783
1279 761
3 5 7 0 0 8320 0 24 31 0 0 3
1270 782
1270 761
1241 761
0 5 8 0 0 8320 0 0 27 187 0 4
964 866
964 857
1352 857
1352 761
0 2 9 0 0 8192 0 0 25 223 0 3
574 857
774 857
774 625
1 2 10 0 0 8320 0 25 26 0 0 3
759 614
759 616
728 616
8 3 11 0 0 4224 0 115 25 0 0 4
1082 584
795 584
795 614
789 614
1 0 12 0 0 8192 0 26 0 0 92 3
692 616
692 605
675 605
0 2 8 0 0 0 0 0 43 187 0 3
606 814
606 604
629 604
0 1 13 0 0 20608 0 0 71 696 0 8
1251 2153
1251 1891
1698 1891
1698 1419
1638 1419
1638 432
1971 432
1971 514
1 0 14 0 0 12416 0 69 0 0 697 8
2183 520
2183 437
1644 437
1644 1424
1694 1424
1694 1898
1241 1898
1241 2105
0 1 15 0 0 20608 0 0 68 698 0 8
1233 2061
1233 1906
1689 1906
1689 1430
1652 1430
1652 443
2481 443
2481 521
1 0 16 0 0 8320 0 67 0 0 699 10
2782 526
2782 451
1658 451
1658 1436
1680 1436
1680 1914
1223 1914
1223 2007
1228 2007
1228 2022
8 0 17 0 0 12288 0 304 0 0 143 5
1206 2259
1215 2259
1215 1922
1672 1922
1672 1536
0 0 9 0 0 8192 0 0 0 277 223 3
250 742
194 742
194 1051
0 2 18 0 0 4096 0 0 46 189 0 3
745 339
745 230
754 230
3 0 19 0 0 4096 0 27 0 0 24 2
1347 716
1347 682
4 0 20 0 0 4096 0 27 0 0 198 2
1338 716
1338 706
2 0 21 0 0 4096 0 27 0 0 73 2
1356 716
1356 643
1 0 22 0 0 4096 0 27 0 0 86 2
1365 716
1365 629
0 0 19 0 0 8320 0 0 0 0 71 4
1386 716
1386 682
907 682
907 664
0 2 23 0 0 8320 0 0 88 0 0 3
1391 717
1391 669
947 669
4 0 24 0 0 4096 0 35 0 0 72 2
1302 716
1302 694
3 0 19 0 0 0 0 35 0 0 24 2
1311 716
1311 682
2 0 21 0 0 0 0 35 0 0 73 2
1320 716
1320 643
1 0 22 0 0 0 0 35 0 0 86 2
1329 716
1329 629
4 0 20 0 0 0 0 30 0 0 198 2
1265 716
1265 706
3 0 23 0 0 0 0 30 0 0 25 2
1274 716
1274 669
2 0 21 0 0 0 0 30 0 0 73 2
1283 716
1283 643
1 0 22 0 0 0 0 30 0 0 86 2
1292 716
1292 629
2 0 21 0 0 0 0 31 0 0 73 2
1245 716
1245 643
3 0 23 0 0 0 0 31 0 0 25 2
1236 716
1236 669
4 0 24 0 0 0 0 31 0 0 72 2
1227 716
1227 694
1 0 22 0 0 0 0 31 0 0 86 2
1254 716
1254 629
4 0 20 0 0 0 0 32 0 0 198 2
1189 716
1189 706
3 0 19 0 0 0 0 32 0 0 24 2
1198 716
1198 682
2 0 25 0 0 4096 0 32 0 0 197 2
1207 716
1207 656
1 0 26 0 0 4096 0 32 0 0 70 2
1216 716
1216 614
3 0 19 0 0 0 0 36 0 0 24 2
1161 716
1161 682
2 0 25 0 0 0 0 36 0 0 197 2
1170 716
1170 656
1 0 26 0 0 0 0 36 0 0 70 2
1179 716
1179 614
4 0 24 0 0 0 0 36 0 0 72 2
1152 716
1152 694
1 0 26 0 0 0 0 33 0 0 70 2
1141 716
1141 614
2 0 25 0 0 0 0 33 0 0 197 2
1132 716
1132 656
3 0 23 0 0 0 0 33 0 0 25 2
1123 716
1123 669
4 0 20 0 0 0 0 33 0 0 198 2
1114 716
1114 706
1 0 26 0 0 0 0 34 0 0 70 2
1105 716
1105 614
2 0 25 0 0 0 0 34 0 0 197 2
1096 716
1096 656
3 0 23 0 0 0 0 34 0 0 25 2
1087 716
1087 669
4 0 24 0 0 0 0 34 0 0 72 2
1078 716
1078 694
1 0 26 0 0 0 0 37 0 0 70 2
1070 716
1070 614
2 0 21 0 0 0 0 37 0 0 73 2
1061 716
1061 643
3 0 19 0 0 0 0 37 0 0 24 2
1052 716
1052 682
4 0 20 0 0 0 0 37 0 0 198 2
1043 716
1043 706
1 0 26 0 0 0 0 39 0 0 70 2
1036 716
1036 614
2 0 21 0 0 0 0 39 0 0 73 2
1027 716
1027 643
3 0 19 0 0 0 0 39 0 0 24 2
1018 716
1018 682
4 0 24 0 0 0 0 39 0 0 72 2
1009 716
1009 694
1 0 26 0 0 0 0 40 0 0 70 2
1001 716
1001 614
2 0 21 0 0 0 0 40 0 0 73 2
992 716
992 643
3 0 23 0 0 0 0 40 0 0 25 2
983 716
983 669
4 0 20 0 0 0 0 40 0 0 198 2
974 716
974 706
1 0 26 0 0 0 0 41 0 0 70 2
966 716
966 614
2 2 21 0 0 0 0 41 87 0 0 3
957 716
955 716
955 643
3 2 23 0 0 0 0 41 88 0 0 3
948 716
947 716
947 669
4 2 24 0 0 0 0 41 113 0 0 3
939 716
938 716
938 694
0 2 26 0 0 8320 0 0 38 0 0 3
1411 719
1411 614
960 614
3 1 19 0 0 0 0 120 88 0 0 4
900 419
907 419
907 669
911 669
0 2 24 0 0 8320 0 0 113 0 0 3
1381 717
1381 694
938 694
0 2 21 0 0 8320 0 0 87 0 0 3
1400 720
1400 643
955 643
0 4 27 0 0 4096 0 0 24 164 0 4
1063 881
1241 881
1241 828
1279 828
1 5 28 0 0 12416 0 28 32 0 0 4
1182 766
1186 766
1186 761
1203 761
2 5 29 0 0 12416 0 28 36 0 0 4
1164 766
1164 764
1166 764
1166 761
0 3 30 0 0 4096 0 0 28 165 0 3
1121 837
1173 837
1173 812
0 3 31 0 0 8192 0 0 29 91 0 4
1026 826
1026 816
1104 816
1104 812
1 5 32 0 0 12416 0 29 33 0 0 4
1113 766
1118 766
1118 761
1128 761
2 5 33 0 0 8320 0 29 34 0 0 3
1095 766
1092 766
1092 761
2 5 34 0 0 8320 0 42 39 0 0 4
990 778
990 768
1023 768
1023 761
1 5 35 0 0 4224 0 42 37 0 0 3
999 778
1057 778
1057 761
3 5 36 0 0 4224 0 42 40 0 0 3
981 778
981 761
988 761
4 5 37 0 0 4224 0 42 41 0 0 3
972 778
953 778
953 761
1 0 22 0 0 0 0 38 0 0 86 2
924 614
923 614
0 3 22 0 0 8320 0 0 44 0 0 5
1406 712
1406 629
923 629
923 212
904 212
1 0 25 0 0 0 0 87 0 0 197 2
919 643
918 643
1 0 20 0 0 0 0 113 0 0 198 2
902 694
901 694
2 5 38 0 0 12416 0 47 42 0 0 5
928 888
915 888
915 832
986 832
986 828
2 0 39 0 0 12416 0 102 0 0 166 5
429 1344
698 1344
698 1264
994 1264
994 1168
0 1 31 0 0 8320 0 0 86 0 0 5
1033 826
1012 826
1012 1228
764 1228
764 1333
9 3 12 0 0 4224 0 48 43 0 0 3
1010 578
675 578
675 613
0 1 40 0 0 8320 0 0 43 274 0 4
275 893
539 893
539 622
629 622
1 13 41 0 0 8320 0 46 115 0 0 5
754 212
754 162
1202 162
1202 539
1146 539
8 1 42 0 0 12416 0 48 115 0 0 4
1034 542
1040 542
1040 521
1082 521
4 0 43 0 0 8320 0 48 0 0 98 3
986 542
846 542
846 212
2 0 9 0 0 0 0 44 0 0 200 3
889 223
915 223
915 332
1 0 43 0 0 0 0 44 0 0 99 2
874 212
809 212
1 4 43 0 0 0 0 45 46 0 0 3
809 201
809 212
802 212
1 0 30 0 0 12288 0 93 0 0 165 4
764 1371
736 1371
736 1241
1032 1241
0 3 3 0 0 12288 0 0 49 228 0 4
656 1588
510 1588
510 1628
280 1628
1 0 44 0 0 12416 0 48 0 0 255 5
986 506
957 506
957 560
866 560
866 519
2 0 45 0 0 16512 0 48 0 0 256 5
986 518
963 518
963 555
859 555
859 419
3 0 46 0 0 16512 0 48 0 0 201 5
986 530
969 530
969 550
852 550
852 321
1 0 44 0 0 0 0 116 0 0 255 2
815 504
815 519
1 0 45 0 0 0 0 119 0 0 256 2
814 404
814 419
1 0 46 0 0 0 0 89 0 0 201 2
813 306
813 321
7 2 47 0 0 4224 0 48 115 0 0 2
1034 530
1082 530
6 3 48 0 0 4224 0 48 115 0 0 4
1034 518
1059 518
1059 539
1082 539
4 5 49 0 0 8320 0 115 48 0 0 4
1082 548
1048 548
1048 506
1034 506
1 0 50 0 0 4224 0 47 0 0 192 2
928 879
414 879
0 2 51 0 0 8320 0 0 49 231 0 5
755 1431
755 1583
504 1583
504 1619
280 1619
2 6 52 0 0 0 0 50 365 0 0 2
379 1787
379 1787
1 3 53 0 0 4224 0 50 51 0 0 4
343 1787
343 1797
344 1797
344 1807
0 9 54 0 0 12416 0 0 52 133 0 5
220 1622
220 1636
170 1636
170 1097
346 1097
3 4 55 0 0 8320 0 134 52 0 0 6
261 421
534 421
534 961
305 961
305 1061
322 1061
3 3 56 0 0 8320 0 131 52 0 0 6
263 516
528 516
528 956
311 956
311 1049
322 1049
3 2 57 0 0 8320 0 125 52 0 0 6
263 606
523 606
523 950
317 950
317 1037
322 1037
3 1 58 0 0 16512 0 128 52 0 0 7
265 701
294 701
294 674
519 674
519 944
322 944
322 1025
8 2 59 0 0 8320 0 54 55 0 0 6
190 1546
175 1546
175 1176
401 1176
401 1145
440 1145
7 2 60 0 0 8320 0 54 56 0 0 6
190 1534
180 1534
180 1183
397 1183
397 1111
440 1111
6 2 61 0 0 8320 0 54 57 0 0 6
190 1522
185 1522
185 1189
393 1189
393 1077
441 1077
5 2 62 0 0 4224 0 54 58 0 0 5
190 1510
190 1195
389 1195
389 1043
442 1043
8 1 63 0 0 8320 0 52 55 0 0 3
370 1061
370 1127
440 1127
7 1 64 0 0 12416 0 52 56 0 0 4
370 1049
376 1049
376 1093
440 1093
6 1 65 0 0 12416 0 52 57 0 0 4
370 1037
384 1037
384 1059
441 1059
5 1 66 0 0 4224 0 52 58 0 0 2
370 1025
442 1025
0 1 67 0 0 4096 0 0 54 224 0 4
759 1545
270 1545
270 1510
238 1510
2 0 68 0 0 12288 0 54 0 0 225 4
238 1522
266 1522
266 1549
747 1549
3 0 69 0 0 12288 0 54 0 0 226 4
238 1534
261 1534
261 1553
735 1553
4 0 70 0 0 12288 0 54 0 0 227 4
238 1546
256 1546
256 1557
723 1557
1 0 71 0 0 12288 0 49 0 0 139 4
280 1610
328 1610
328 1579
479 1579
1 4 54 0 0 0 0 53 49 0 0 4
214 1622
226 1622
226 1619
235 1619
2 9 72 0 0 4224 0 53 54 0 0 2
214 1586
214 1582
3 4 73 0 0 8320 0 55 535 0 0 4
486 1136
495 1136
495 1092
503 1092
3 3 74 0 0 8320 0 56 535 0 0 4
486 1102
491 1102
491 1080
503 1080
3 2 75 0 0 4224 0 57 535 0 0 2
487 1068
503 1068
3 1 76 0 0 8320 0 58 535 0 0 4
488 1034
491 1034
491 1056
503 1056
0 1 71 0 0 12416 0 0 59 782 0 5
479 1697
479 1564
622 1564
622 1396
644 1396
0 5 39 0 0 0 0 0 47 166 0 4
1001 900
993 900
993 892
978 892
0 3 77 0 0 4224 0 0 306 244 0 4
707 1910
707 2344
1043 2344
1043 2332
0 1 17 0 0 0 0 0 65 143 0 3
1674 634
1674 635
1678 635
3 1 17 0 0 8320 0 60 70 0 0 7
1656 1536
1674 1536
1674 471
1816 471
1816 537
1824 537
1824 582
2 0 3 0 0 12416 0 60 0 0 228 4
1611 1545
1582 1545
1582 1520
815 1520
0 1 78 0 0 4224 0 0 60 344 0 4
632 1512
1593 1512
1593 1527
1611 1527
0 0 79 0 0 16384 0 0 0 147 158 5
1905 516
1905 544
1873 544
1873 635
1754 635
2 2 79 0 0 0 0 64 63 0 0 8
1894 510
1894 516
1932 516
1932 507
2034 507
2034 519
2116 519
2116 510
0 2 79 0 0 12288 0 0 63 149 0 5
2432 505
2411 505
2411 513
2116 513
2116 510
2 2 79 0 0 8320 0 61 62 0 0 4
2731 493
2731 505
2432 505
2432 498
2 3 80 0 0 4224 0 67 61 0 0 3
2764 526
2764 482
2746 482
2 3 81 0 0 4224 0 68 62 0 0 3
2463 521
2463 487
2447 487
2 3 82 0 0 8320 0 69 63 0 0 3
2165 520
2165 499
2131 499
1 1 83 0 0 4224 0 61 2 0 0 2
2716 482
2711 482
1 1 84 0 0 4224 0 62 3 0 0 2
2417 487
2412 487
1 1 85 0 0 4224 0 63 4 0 0 2
2101 499
2096 499
3 2 86 0 0 4224 0 64 71 0 0 3
1909 499
1953 499
1953 514
1 1 87 0 0 4224 0 64 5 0 0 2
1879 499
1874 499
2 2 79 0 0 0 0 66 65 0 0 5
1754 569
1754 567
1754 567
1754 635
1714 635
2 3 88 0 0 8320 0 70 66 0 0 3
1806 582
1806 558
1769 558
1 1 89 0 0 4224 0 66 6 0 0 2
1739 558
1734 558
3 0 90 0 0 0 0 70 0 0 1174 2
1815 628
1815 628
1 3 91 0 0 8320 0 530 67 0 0 3
2783 590
2773 590
2773 572
3 0 92 0 0 4224 0 47 0 0 772 3
928 897
640 897
640 1009
1 0 27 0 0 16512 0 92 0 0 0 7
764 1413
743 1413
743 1233
1017 1233
1017 937
1063 937
1063 871
0 2 30 0 0 12416 0 0 79 0 0 7
1125 833
1125 837
1032 837
1032 1402
1271 1402
1271 1396
1310 1396
2 1 39 0 0 0 0 81 77 0 0 5
970 1168
1001 1168
1001 893
1128 893
1128 898
1 8 93 0 0 8320 0 103 76 0 0 4
1186 1184
1159 1184
1159 965
1152 965
7 1 94 0 0 8320 0 76 104 0 0 4
1152 977
1166 977
1166 1153
1188 1153
1 6 95 0 0 8320 0 105 76 0 0 4
1189 1122
1174 1122
1174 989
1152 989
1 5 96 0 0 8320 0 106 76 0 0 4
1191 1091
1182 1091
1182 1001
1152 1001
0 4 97 0 0 4096 0 0 76 245 0 3
1072 1095
1072 965
1104 965
0 3 98 0 0 4096 0 0 76 246 0 3
1064 1080
1064 977
1104 977
0 2 99 0 0 4096 0 0 76 247 0 3
1057 1069
1057 989
1104 989
1 0 100 0 0 4096 0 76 0 0 248 3
1104 1001
1049 1001
1049 1056
2 9 101 0 0 4224 0 77 76 0 0 2
1128 934
1128 929
0 0 102 0 0 8192 0 0 0 784 341 3
504 1715
504 1711
495 1711
1 0 31 0 0 0 0 78 0 0 91 4
875 1358
868 1358
868 1309
764 1309
9 2 103 0 0 8320 0 80 78 0 0 7
1224 1387
1224 1395
971 1395
971 1367
923 1367
923 1358
911 1358
1 10 104 0 0 8320 0 80 154 0 0 4
1200 1315
1174 1315
1174 1352
1164 1352
2 11 105 0 0 12416 0 80 154 0 0 4
1200 1327
1194 1327
1194 1343
1164 1343
3 12 106 0 0 4224 0 80 154 0 0 4
1200 1339
1180 1339
1180 1334
1164 1334
13 4 107 0 0 8320 0 154 80 0 0 4
1164 1325
1186 1325
1186 1351
1200 1351
2 8 108 0 0 12416 0 103 80 0 0 6
1187 1193
1112 1193
1112 1237
1275 1237
1275 1351
1248 1351
7 2 109 0 0 12416 0 80 104 0 0 6
1248 1339
1269 1339
1269 1244
1105 1244
1105 1162
1189 1162
6 2 110 0 0 12416 0 80 105 0 0 6
1248 1327
1257 1327
1257 1253
1098 1253
1098 1131
1190 1131
5 2 111 0 0 12416 0 80 106 0 0 5
1248 1315
1248 1268
1092 1268
1092 1100
1192 1100
1 0 8 0 0 0 0 83 0 0 0 4
589 814
921 814
921 866
974 866
3 9 112 0 0 4224 0 81 82 0 0 2
959 1153
959 1122
2 2 18 0 0 0 0 91 121 0 0 4
756 339
744 339
744 437
751 437
3 0 113 0 0 4224 0 83 0 0 191 4
559 814
426 814
426 815
425 815
2 2 113 0 0 0 0 85 84 0 0 5
392 836
399 836
399 809
425 809
425 837
0 1 50 0 0 0 0 0 84 257 0 3
296 914
414 914
414 852
2 1 114 0 0 8320 0 122 85 0 0 3
360 899
381 899
381 851
8 3 115 0 0 8320 0 136 84 0 0 4
401 767
387 767
387 822
414 822
3 7 116 0 0 4224 0 85 136 0 0 3
381 821
381 758
401 758
3 8 117 0 0 12416 0 86 154 0 0 6
809 1342
839 1342
839 1420
1057 1420
1057 1370
1100 1370
3 0 25 0 0 12416 0 90 0 0 0 5
905 321
918 321
918 656
1396 656
1396 714
0 3 20 0 0 8320 0 0 117 0 0 5
1377 717
1377 706
901 706
901 519
903 519
12 1 118 0 0 12416 0 115 91 0 0 6
1146 548
1208 548
1208 157
718 157
718 321
756 321
2 0 9 0 0 0 0 90 0 0 252 3
890 332
915 332
915 453
4 1 46 0 0 0 0 91 90 0 0 2
804 321
875 321
3 0 3 0 0 0 0 92 0 0 228 2
809 1422
815 1422
2 0 51 0 0 0 0 93 0 0 231 2
764 1389
755 1389
0 0 9 0 0 4096 0 0 0 222 289 5
823 844
1419 844
1419 675
1806 675
1806 667
1 0 119 0 0 12416 0 97 0 0 218 4
1201 928
1201 959
1249 959
1249 1193
0 1 120 0 0 4224 0 0 96 217 0 4
1255 1162
1255 948
1223 948
1223 928
1 0 121 0 0 8320 0 95 0 0 219 3
1245 928
1259 928
1259 1131
1 0 122 0 0 4224 0 94 0 0 220 2
1268 928
1268 1100
1 0 123 0 0 4096 0 101 0 0 1102 2
892 955
892 1092
1 0 124 0 0 4096 0 100 0 0 1103 2
908 955
908 1080
0 1 125 0 0 12288 0 0 99 1104 0 4
918 1068
918 1030
924 1030
924 955
0 1 126 0 0 12288 0 0 98 1105 0 4
922 1056
922 1034
940 1034
940 955
5 3 127 0 0 8320 0 110 106 0 0 5
1425 1287
1425 1227
1127 1227
1127 1109
1191 1109
6 3 128 0 0 8320 0 110 105 0 0 5
1413 1287
1413 1223
1133 1223
1133 1140
1189 1140
7 3 129 0 0 8320 0 110 104 0 0 5
1401 1287
1401 1218
1138 1218
1138 1171
1188 1171
8 3 130 0 0 8320 0 110 103 0 0 5
1389 1287
1389 1213
1142 1213
1142 1202
1186 1202
2 4 120 0 0 0 0 538 104 0 0 4
1313 1128
1302 1128
1302 1162
1234 1162
1 4 119 0 0 0 0 538 103 0 0 4
1313 1137
1310 1137
1310 1193
1232 1193
3 4 121 0 0 0 0 538 105 0 0 4
1313 1119
1295 1119
1295 1131
1235 1131
4 4 122 0 0 0 0 106 538 0 0 4
1237 1100
1299 1100
1299 1110
1313 1110
1 0 9 0 0 12416 0 51 0 0 289 4
298 1798
291 1798
291 1502
1855 1502
0 0 9 0 0 0 0 0 0 0 223 6
838 692
823 692
823 928
287 928
287 1051
280 1051
1 2 9 0 0 0 0 1 83 0 0 5
146 1051
281 1051
281 921
574 921
574 825
1 0 67 0 0 0 0 155 0 0 806 2
759 1799
759 1485
2 0 68 0 0 0 0 155 0 0 807 2
747 1799
747 1473
3 0 69 0 0 0 0 155 0 0 808 2
735 1799
735 1461
4 0 70 0 0 0 0 155 0 0 809 2
723 1799
723 1449
1 0 3 0 0 0 0 111 0 0 202 5
656 1901
656 1520
815 1520
815 1422
812 1422
2 0 51 0 0 0 0 107 0 0 231 2
748 1424
755 1424
4 1 50 0 0 0 0 59 107 0 0 4
696 1405
707 1405
707 1424
712 1424
2 2 51 0 0 0 0 86 92 0 0 4
764 1351
755 1351
755 1431
764 1431
1 0 67 0 0 0 0 109 0 0 806 2
1425 1395
1425 1485
2 0 68 0 0 0 0 109 0 0 807 2
1413 1395
1413 1473
3 0 69 0 0 0 0 109 0 0 808 2
1401 1395
1401 1461
4 0 70 0 0 0 0 109 0 0 809 2
1389 1395
1389 1449
2 9 131 0 0 0 0 108 110 0 0 2
1353 1311
1353 1311
0 1 132 0 0 8192 0 0 79 1182 0 4
959 1301
959 1408
1295 1408
1295 1407
3 9 133 0 0 4224 0 79 109 0 0 3
1325 1407
1325 1371
1359 1371
4 8 134 0 0 4224 0 110 109 0 0 2
1389 1335
1389 1347
3 7 135 0 0 4224 0 110 109 0 0 2
1401 1335
1401 1347
2 6 136 0 0 4224 0 110 109 0 0 2
1413 1335
1413 1347
1 5 137 0 0 4224 0 110 109 0 0 2
1425 1335
1425 1347
9 2 138 0 0 8320 0 155 112 0 0 4
687 1823
687 1869
750 1869
750 1910
1 3 77 0 0 0 0 112 111 0 0 2
714 1910
701 1910
8 1 97 0 0 8320 0 82 154 0 0 4
983 1092
1072 1092
1072 1307
1100 1307
7 2 98 0 0 8320 0 82 154 0 0 4
983 1080
1064 1080
1064 1316
1100 1316
3 6 99 0 0 8320 0 154 82 0 0 4
1100 1325
1057 1325
1057 1068
983 1068
5 4 100 0 0 8320 0 82 154 0 0 4
983 1056
1049 1056
1049 1334
1100 1334
3 0 18 0 0 8320 0 114 0 0 250 3
695 714
744 714
744 537
2 2 18 0 0 0 0 121 118 0 0 4
751 437
744 437
744 537
754 537
0 0 9 0 0 0 0 0 0 252 222 4
888 540
888 605
825 605
825 692
2 2 9 0 0 0 0 120 117 0 0 6
885 430
885 453
915 453
915 540
888 540
888 530
1 11 139 0 0 12416 0 121 115 0 0 6
751 419
713 419
713 147
1215 147
1215 557
1146 557
10 1 140 0 0 12416 0 115 118 0 0 6
1146 566
1224 566
1224 133
707 133
707 519
754 519
4 1 44 0 0 0 0 118 117 0 0 2
802 519
873 519
4 1 45 0 0 0 0 121 120 0 0 2
799 419
870 419
0 1 50 0 0 0 0 0 122 230 0 7
704 1405
704 1404
707 1404
707 1206
296 1206
296 899
324 899
3 0 141 0 0 8320 0 123 0 0 283 3
252 836
210 836
210 516
0 0 132 0 0 8320 0 0 0 262 1183 5
107 719
17 719
17 1213
431 1213
431 1301
2 0 132 0 0 0 0 130 0 0 262 2
114 534
107 534
2 0 132 0 0 0 0 124 0 0 262 2
114 624
107 624
2 2 132 0 0 0 0 135 129 0 0 4
112 439
107 439
107 719
116 719
1 10 142 0 0 12416 0 129 136 0 0 6
116 701
90 701
90 368
499 368
499 749
465 749
1 11 143 0 0 12416 0 124 136 0 0 6
114 606
95 606
95 360
490 360
490 740
465 740
1 12 144 0 0 12416 0 130 136 0 0 6
114 516
102 516
102 351
482 351
482 731
465 731
1 13 145 0 0 12416 0 135 136 0 0 5
112 421
112 343
474 343
474 722
465 722
4 0 146 0 0 8320 0 123 0 0 285 3
252 848
204 848
204 421
2 0 147 0 0 8320 0 123 0 0 281 3
252 824
218 824
218 606
1 0 148 0 0 8320 0 123 0 0 279 3
252 812
226 812
226 701
8 1 149 0 0 8320 0 123 136 0 0 4
300 848
330 848
330 704
401 704
7 2 150 0 0 8320 0 123 136 0 0 4
300 836
340 836
340 713
401 713
6 3 151 0 0 8320 0 123 136 0 0 4
300 824
350 824
350 722
401 722
5 4 152 0 0 8320 0 123 136 0 0 4
300 812
360 812
360 731
401 731
1 9 40 0 0 0 0 8 123 0 0 3
231 893
276 893
276 884
2 0 9 0 0 0 0 131 0 0 277 2
248 527
301 527
2 0 9 0 0 0 0 125 0 0 277 2
248 617
301 617
2 2 9 0 0 0 0 134 128 0 0 6
246 432
246 446
301 446
301 742
250 742
250 712
1 0 148 0 0 0 0 127 0 0 279 2
195 686
195 701
4 1 148 0 0 0 0 129 128 0 0 2
164 701
235 701
1 0 147 0 0 0 0 126 0 0 281 2
193 591
193 606
4 1 147 0 0 0 0 124 125 0 0 2
162 606
233 606
1 0 141 0 0 0 0 132 0 0 283 2
193 501
193 516
4 1 141 0 0 0 0 130 131 0 0 2
162 516
233 516
1 0 146 0 0 0 0 133 0 0 285 2
191 406
191 421
4 1 146 0 0 0 0 135 134 0 0 2
160 421
231 421
0 0 153 0 0 8192 0 0 0 810 945 4
1824 1662
1824 1678
1870 1678
1870 1662
3 9 154 0 0 4224 0 137 375 0 0 2
3080 1697
3080 1693
1 0 153 0 0 0 0 137 0 0 945 2
3080 1667
3080 1661
0 2 9 0 0 0 0 0 137 0 0 10
1788 667
1855 667
1855 1645
1843 1645
1843 1650
1954 1650
1954 1668
3060 1668
3060 1682
3069 1682
5 1 155 0 0 8320 0 538 22 0 0 3
1313 1083
1285 1083
1285 1037
6 1 156 0 0 8320 0 538 21 0 0 3
1307 1065
1306 1065
1306 1037
0 1 90 0 0 4096 0 0 138 304 0 3
3089 1258
3089 1490
3078 1490
0 1 157 0 0 12288 0 0 418 911 0 4
3078 1460
3116 1460
3116 1521
3050 1521
2 3 158 0 0 8320 0 402 138 0 0 3
3031 1458
3033 1458
3033 1481
0 1 90 0 0 4096 0 0 139 307 0 3
2771 1257
2771 1494
2750 1494
1 0 159 0 0 8192 0 424 0 0 912 4
2724 1525
2794 1525
2794 1454
2750 1454
2 3 160 0 0 8320 0 403 139 0 0 3
2706 1460
2705 1460
2705 1485
0 1 90 0 0 0 0 0 140 310 0 3
2487 1259
2487 1489
2462 1489
1 0 161 0 0 8192 0 430 0 0 913 4
2436 1523
2495 1523
2495 1456
2462 1456
2 3 162 0 0 8320 0 404 140 0 0 3
2415 1460
2417 1460
2417 1480
0 1 90 0 0 0 0 0 141 313 0 3
2194 1263
2194 1493
2173 1493
1 0 163 0 0 8192 0 436 0 0 914 4
2145 1526
2206 1526
2206 1460
2173 1460
2 3 164 0 0 4224 0 405 141 0 0 3
2122 1461
2122 1484
2128 1484
0 1 90 0 0 0 0 0 142 316 0 6
3074 1037
3079 1037
3079 1181
3089 1181
3089 1259
3082 1259
1 0 165 0 0 8192 0 442 0 0 915 4
3056 1288
3103 1288
3103 1230
3083 1230
3 2 166 0 0 8320 0 142 398 0 0 3
3037 1250
3036 1250
3036 1226
0 1 90 0 0 0 0 0 143 319 0 3
2771 1046
2771 1258
2759 1258
0 1 167 0 0 12288 0 0 448 916 0 4
2760 1231
2792 1231
2792 1290
2730 1290
3 2 168 0 0 8320 0 143 399 0 0 4
2714 1249
2706 1249
2706 1227
2711 1227
0 1 90 0 0 0 0 0 144 323 0 3
2487 1038
2487 1259
2473 1259
1 0 169 0 0 8192 0 454 0 0 917 4
2442 1287
2493 1287
2493 1218
2474 1218
3 2 170 0 0 4224 0 144 400 0 0 3
2428 1250
2428 1224
2424 1224
1 0 90 0 0 0 0 145 0 0 326 3
2183 1263
2195 1263
2195 1041
1 0 171 0 0 8192 0 460 0 0 918 4
2151 1290
2205 1290
2205 1227
2183 1227
2 3 172 0 0 4224 0 401 145 0 0 3
2132 1226
2132 1254
2138 1254
0 1 90 0 0 0 0 0 146 329 0 5
3078 820
3078 842
3074 842
3074 1042
3071 1042
1 0 173 0 0 8192 0 466 0 0 919 4
3059 1072
3088 1072
3088 1010
3081 1010
3 2 174 0 0 4224 0 146 406 0 0 3
3026 1033
3026 1010
3038 1010
1 0 90 0 0 0 0 147 0 0 320 3
2755 1046
2771 1046
2771 821
1 0 90 0 0 0 0 151 0 0 1174 3
2761 821
2771 821
2771 628
1 0 175 0 0 8192 0 472 0 0 920 4
2733 1075
2793 1075
2793 1010
2755 1010
2 3 176 0 0 4224 0 407 147 0 0 2
2710 1010
2710 1037
0 1 90 0 0 0 0 0 148 336 0 3
2487 821
2487 1038
2471 1038
1 0 177 0 0 8192 0 478 0 0 921 4
2445 1070
2493 1070
2493 1003
2475 1003
2 3 178 0 0 4224 0 408 148 0 0 2
2426 1007
2426 1029
1 0 90 0 0 0 0 149 0 0 334 3
2185 1046
2195 1046
2195 823
1 0 179 0 0 8192 0 484 0 0 922 4
2154 1075
2205 1075
2205 1013
2186 1013
2 3 180 0 0 4224 0 409 149 0 0 3
2136 1010
2136 1037
2140 1037
1 0 90 0 0 12288 0 150 0 0 1174 4
3072 820
3079 820
3079 628
2793 628
0 1 181 0 0 8192 0 0 490 923 0 4
3076 789
3083 789
3083 848
3049 848
3 2 182 0 0 8320 0 150 410 0 0 3
3027 811
3025 811
3025 788
0 1 183 0 0 8192 0 0 496 924 0 4
2761 788
2785 788
2785 854
2735 854
3 2 184 0 0 4224 0 151 411 0 0 2
2716 812
2716 790
1 0 90 0 0 0 0 153 0 0 1174 5
2190 823
2195 823
2195 645
2188 645
2188 628
2 0 185 0 0 4096 0 153 0 0 340 2
2190 805
2203 805
1 0 90 0 0 0 0 152 0 0 1174 3
2479 821
2487 821
2487 628
1 0 186 0 0 8192 0 502 0 0 925 4
2454 850
2493 850
2493 785
2479 785
3 2 187 0 0 8320 0 152 412 0 0 3
2434 812
2435 812
2435 789
2 3 188 0 0 4224 0 509 153 0 0 3
2137 794
2137 814
2145 814
0 1 185 0 0 8320 0 0 508 1184 0 7
1446 926
1446 789
1915 789
1915 707
2203 707
2203 856
2153 856
3 2 102 0 0 12416 0 59 111 0 0 7
644 1414
644 1578
495 1578
495 1918
624 1918
624 1919
656 1919
9 3 189 0 0 8320 0 536 102 0 0 4
579 1419
579 1389
418 1389
418 1359
1 0 132 0 0 0 0 102 0 0 1182 4
418 1329
418 1312
585 1312
585 1301
0 2 78 0 0 0 0 0 59 783 0 5
487 1706
487 1571
632 1571
632 1405
645 1405
2 8 190 0 0 16512 0 75 155 0 0 6
931 1972
931 1907
925 1907
925 1860
723 1860
723 1847
2 7 191 0 0 16512 0 74 155 0 0 6
971 1974
971 1908
966 1908
966 1855
735 1855
735 1847
2 6 192 0 0 12416 0 73 155 0 0 5
1007 1973
1005 1973
1005 1851
747 1851
747 1847
2 5 193 0 0 8320 0 72 155 0 0 3
1044 1971
1044 1847
759 1847
1 8 194 0 0 16512 0 75 345 0 0 6
940 1971
940 1908
943 1908
943 1859
1062 1859
1062 1832
1 7 195 0 0 16512 0 74 345 0 0 6
980 1973
980 1910
984 1910
984 1863
1074 1863
1074 1832
1 6 196 0 0 4224 0 73 345 0 0 6
1016 1972
1016 1883
1023 1883
1023 1867
1086 1867
1086 1832
1 5 197 0 0 4224 0 72 345 0 0 6
1053 1970
1053 1885
1062 1885
1062 1871
1098 1871
1098 1832
7 0 198 0 0 12288 0 302 0 0 384 4
1887 2268
1887 2509
1552 2509
1552 3139
3 8 199 0 0 4224 0 156 303 0 0 4
1256 2874
1256 2506
1547 2506
1547 2263
2 0 198 0 0 0 0 156 0 0 384 2
1265 2920
1265 3139
1 0 200 0 0 4096 0 156 0 0 393 2
1247 2920
1247 2954
7 0 200 0 0 4096 0 304 0 0 393 2
1197 2259
1197 2954
6 0 201 0 0 16384 0 302 0 0 394 6
1878 2268
1878 2341
1883 2341
1883 2501
1546 2501
1546 2757
7 0 201 0 0 4096 0 303 0 0 394 2
1538 2263
1538 2757
0 2 202 0 0 16512 0 0 256 414 0 6
1976 3226
2077 3226
2077 2933
2725 2933
2725 1990
2737 1990
0 2 203 0 0 16512 0 0 248 415 0 6
1963 3214
2072 3214
2072 2927
2719 2927
2719 2116
2735 2116
0 2 204 0 0 16512 0 0 244 416 0 6
1950 3202
2067 3202
2067 2923
2714 2923
2714 2238
2734 2238
0 2 205 0 0 12416 0 0 240 417 0 6
1937 3190
2059 3190
2059 2917
2709 2917
2709 2361
2734 2361
0 1 206 0 0 16512 0 0 256 423 0 6
1976 3041
2051 3041
2051 2910
2704 2910
2704 1972
2737 1972
0 1 207 0 0 16512 0 0 248 424 0 6
1963 3029
2041 3029
2041 2903
2699 2903
2699 2098
2735 2098
0 1 208 0 0 16512 0 0 244 425 0 6
1950 3016
2034 3016
2034 2895
2695 2895
2695 2220
2734 2220
1 0 209 0 0 12416 0 240 0 0 426 6
2734 2343
2692 2343
2692 2889
2028 2889
2028 3005
1933 3005
0 1 210 0 0 16512 0 0 254 432 0 6
1973 2844
2030 2844
2030 2884
2689 2884
2689 1958
2735 1958
0 1 211 0 0 16512 0 0 250 433 0 6
1958 2832
2036 2832
2036 2879
2684 2879
2684 2078
2734 2078
0 1 212 0 0 16512 0 0 246 434 0 6
1947 2819
2040 2819
2040 2874
2681 2874
2681 2203
2733 2203
0 1 213 0 0 12416 0 0 242 435 0 6
1933 2808
2044 2808
2044 2870
2675 2870
2675 2325
2732 2325
0 2 214 0 0 16512 0 0 254 441 0 6
1971 2663
2050 2663
2050 2865
2671 2865
2671 1949
2735 1949
0 2 215 0 0 16512 0 0 250 442 0 6
1959 2651
2055 2651
2055 2860
2666 2860
2666 2069
2734 2069
0 2 216 0 0 16512 0 0 246 443 0 6
1946 2639
2060 2639
2060 2855
2661 2855
2661 2194
2733 2194
0 2 217 0 0 12416 0 0 242 444 0 6
1933 2627
2064 2627
2064 2851
2657 2851
2657 2316
2732 2316
0 2 218 0 0 4096 0 0 166 395 0 3
1604 2892
1604 3275
1679 3275
0 2 219 0 0 4096 0 0 165 396 0 3
1614 2859
1614 3240
1680 3240
0 2 220 0 0 4096 0 0 164 397 0 3
1624 2824
1624 3206
1680 3206
0 2 221 0 0 4096 0 0 163 398 0 3
1636 2791
1636 3173
1680 3173
1 0 222 0 0 8192 0 166 0 0 385 3
1679 3257
1562 3257
1562 3090
0 1 223 0 0 4096 0 0 165 386 0 3
1568 3055
1568 3222
1680 3222
0 1 224 0 0 4096 0 0 164 387 0 3
1575 3021
1575 3188
1680 3188
1 0 225 0 0 8192 0 163 0 0 388 3
1680 3155
1580 3155
1580 2988
0 1 198 0 0 4224 0 0 158 785 0 5
502 1724
502 2523
1069 2523
1069 3139
1856 3139
2 0 222 0 0 8192 0 167 0 0 399 3
1679 3090
1562 3090
1562 2875
2 0 223 0 0 8192 0 168 0 0 400 3
1680 3055
1568 3055
1568 2841
2 0 224 0 0 8192 0 169 0 0 401 3
1680 3021
1575 3021
1575 2806
2 0 225 0 0 8192 0 170 0 0 402 3
1680 2988
1580 2988
1580 2773
1 0 16 0 0 0 0 167 0 0 407 3
1679 3072
1323 3072
1323 2694
1 0 15 0 0 0 0 168 0 0 408 3
1680 3037
1357 3037
1357 2660
1 0 14 0 0 0 0 169 0 0 409 3
1680 3003
1382 3003
1382 2625
1 0 13 0 0 0 0 170 0 0 410 3
1680 2970
1408 2970
1408 2592
0 1 200 0 0 4224 0 0 175 786 0 5
508 1733
508 2514
1078 2514
1078 2954
1856 2954
0 1 201 0 0 16512 0 0 182 787 0 5
514 1742
514 2503
1087 2503
1087 2757
1853 2757
0 2 218 0 0 0 0 0 180 597 0 5
1907 2194
1907 2532
1604 2532
1604 2893
1681 2893
0 2 219 0 0 0 0 0 179 634 0 5
1914 2182
1914 2538
1614 2538
1614 2859
1681 2859
0 2 220 0 0 0 0 0 178 598 0 5
1919 2170
1919 2547
1624 2547
1624 2824
1681 2824
0 2 221 0 0 4096 0 0 177 633 0 5
1925 2158
1925 2555
1636 2555
1636 2791
1681 2791
0 1 222 0 0 0 0 0 180 403 0 3
1562 2712
1562 2875
1681 2875
0 1 223 0 0 0 0 0 179 404 0 3
1568 2678
1568 2841
1681 2841
1 0 224 0 0 0 0 178 0 0 405 3
1681 2806
1574 2806
1574 2643
1 0 225 0 0 0 0 177 0 0 406 3
1681 2773
1580 2773
1580 2610
0 2 222 0 0 4096 0 0 217 603 0 3
1562 2425
1562 2712
1680 2712
0 2 223 0 0 4096 0 0 218 636 0 3
1568 2431
1568 2678
1680 2678
0 2 224 0 0 0 0 0 219 604 0 3
1574 2437
1574 2643
1680 2643
2 0 225 0 0 0 0 220 0 0 635 3
1680 2610
1580 2610
1580 2443
0 1 16 0 0 0 0 0 217 639 0 3
1285 2399
1285 2694
1680 2694
0 1 15 0 0 0 0 0 218 605 0 3
1293 2406
1293 2660
1680 2660
0 1 14 0 0 0 0 0 219 638 0 3
1302 2413
1302 2625
1680 2625
0 1 13 0 0 0 0 0 220 637 0 3
1311 2420
1311 2592
1680 2592
6 0 226 0 0 4096 0 303 0 0 413 2
1529 2263
1529 2495
6 0 226 0 0 4096 0 304 0 0 413 2
1188 2259
1188 2495
0 1 226 0 0 8320 0 0 191 788 0 5
520 1751
520 2495
1814 2495
1814 2576
1852 2576
5 1 202 0 0 0 0 157 162 0 0 3
1918 3226
1976 3226
1976 3180
6 1 203 0 0 0 0 157 161 0 0 3
1918 3214
1963 3214
1963 3180
1 7 204 0 0 0 0 160 157 0 0 3
1950 3179
1950 3202
1918 3202
8 1 205 0 0 0 0 157 159 0 0 3
1918 3190
1937 3190
1937 3179
3 1 227 0 0 4224 0 166 157 0 0 4
1728 3266
1821 3266
1821 3226
1870 3226
2 3 228 0 0 12416 0 157 165 0 0 4
1870 3214
1804 3214
1804 3231
1729 3231
3 3 229 0 0 4224 0 164 157 0 0 4
1729 3197
1821 3197
1821 3202
1870 3202
4 3 230 0 0 12416 0 157 163 0 0 4
1870 3190
1840 3190
1840 3164
1729 3164
2 9 231 0 0 8320 0 158 157 0 0 3
1892 3139
1894 3139
1894 3154
5 1 206 0 0 0 0 176 171 0 0 3
1918 3041
1976 3041
1976 2995
6 1 207 0 0 0 0 176 172 0 0 3
1918 3029
1963 3029
1963 2995
1 7 208 0 0 0 0 173 176 0 0 3
1950 2994
1950 3017
1918 3017
8 1 209 0 0 0 0 176 174 0 0 3
1918 3005
1937 3005
1937 2994
3 1 232 0 0 4224 0 167 176 0 0 4
1728 3081
1821 3081
1821 3041
1870 3041
2 3 233 0 0 12416 0 176 168 0 0 4
1870 3029
1804 3029
1804 3046
1729 3046
3 3 234 0 0 4224 0 169 176 0 0 4
1729 3012
1821 3012
1821 3017
1870 3017
4 3 235 0 0 12416 0 176 170 0 0 4
1870 3005
1840 3005
1840 2979
1729 2979
2 9 236 0 0 8320 0 175 176 0 0 3
1892 2954
1894 2954
1894 2969
5 1 210 0 0 0 0 181 186 0 0 3
1915 2844
1973 2844
1973 2798
6 1 211 0 0 0 0 181 185 0 0 3
1915 2832
1960 2832
1960 2798
1 7 212 0 0 0 0 184 181 0 0 3
1947 2797
1947 2820
1915 2820
8 1 213 0 0 0 0 181 183 0 0 3
1915 2808
1934 2808
1934 2797
3 1 237 0 0 4224 0 180 181 0 0 4
1727 2884
1818 2884
1818 2844
1867 2844
2 3 238 0 0 12416 0 181 179 0 0 4
1867 2832
1801 2832
1801 2850
1727 2850
3 3 239 0 0 4224 0 178 181 0 0 4
1727 2815
1818 2815
1818 2820
1867 2820
4 3 240 0 0 12416 0 181 177 0 0 4
1867 2808
1837 2808
1837 2782
1727 2782
2 9 241 0 0 8320 0 182 181 0 0 3
1889 2757
1891 2757
1891 2772
5 1 214 0 0 0 0 192 187 0 0 3
1914 2663
1972 2663
1972 2617
6 1 215 0 0 0 0 192 188 0 0 3
1914 2651
1959 2651
1959 2617
1 7 216 0 0 0 0 189 192 0 0 3
1946 2616
1946 2639
1914 2639
8 1 217 0 0 0 0 192 190 0 0 3
1914 2627
1933 2627
1933 2616
3 1 242 0 0 4224 0 217 192 0 0 4
1726 2703
1817 2703
1817 2663
1866 2663
2 3 243 0 0 12416 0 192 218 0 0 4
1866 2651
1800 2651
1800 2669
1726 2669
3 3 244 0 0 4224 0 219 192 0 0 4
1726 2634
1817 2634
1817 2639
1866 2639
4 3 245 0 0 12416 0 192 220 0 0 4
1866 2627
1836 2627
1836 2601
1726 2601
2 9 246 0 0 8320 0 191 192 0 0 3
1888 2576
1890 2576
1890 2591
0 3 247 0 0 8320 0 0 254 473 0 4
2540 2783
2651 2783
2651 1940
2735 1940
0 3 248 0 0 8320 0 0 250 474 0 4
2526 2771
2644 2771
2644 2060
2734 2060
0 3 249 0 0 8320 0 0 246 475 0 4
2516 2757
2638 2757
2638 2185
2733 2185
0 3 250 0 0 8320 0 0 242 476 0 4
2502 2747
2634 2747
2634 2307
2732 2307
0 4 251 0 0 8320 0 0 254 477 0 4
2539 2605
2628 2605
2628 1931
2735 1931
0 4 252 0 0 8320 0 0 250 478 0 4
2525 2593
2623 2593
2623 2051
2734 2051
0 4 253 0 0 8320 0 0 246 479 0 4
2513 2580
2617 2580
2617 2176
2733 2176
0 4 254 0 0 8320 0 0 242 480 0 4
2499 2569
2611 2569
2611 2298
2732 2298
5 0 255 0 0 4096 0 302 0 0 460 2
1869 2268
1869 2525
5 0 255 0 0 0 0 304 0 0 460 2
1179 2259
1179 2486
0 1 255 0 0 8320 0 0 210 789 0 7
527 1760
527 2486
1819 2486
1819 2525
2069 2525
2069 2696
2421 2696
0 2 16 0 0 0 0 0 208 510 0 3
2075 2439
2075 2831
2250 2831
0 2 15 0 0 0 0 0 209 511 0 3
2081 2405
2081 2797
2249 2797
0 2 14 0 0 0 0 0 207 512 0 3
2088 2372
2088 2764
2248 2764
0 2 13 0 0 0 0 0 206 513 0 3
2095 2338
2095 2730
2248 2730
1 0 218 0 0 0 0 208 0 0 469 3
2250 2813
2161 2813
2161 2653
0 1 219 0 0 0 0 0 209 470 0 3
2174 2619
2174 2779
2249 2779
0 1 220 0 0 0 0 0 207 471 0 3
2185 2586
2185 2746
2248 2746
0 1 221 0 0 0 0 0 206 472 0 3
2191 2552
2191 2712
2248 2712
0 2 218 0 0 4096 0 0 214 597 0 3
2104 2194
2104 2653
2247 2653
2 0 219 0 0 8192 0 215 0 0 634 3
2246 2619
2114 2619
2114 2182
0 2 220 0 0 4096 0 0 213 598 0 3
2123 2170
2123 2586
2246 2586
0 2 221 0 0 0 0 0 212 633 0 3
2132 2158
2132 2552
2245 2552
5 1 247 0 0 0 0 205 196 0 0 3
2483 2783
2542 2783
2542 2737
6 1 248 0 0 0 0 205 195 0 0 3
2483 2771
2529 2771
2529 2737
1 7 249 0 0 0 0 194 205 0 0 3
2516 2736
2516 2759
2483 2759
8 1 250 0 0 0 0 205 193 0 0 3
2483 2747
2503 2747
2503 2736
5 1 251 0 0 0 0 211 200 0 0 3
2480 2605
2539 2605
2539 2559
6 1 252 0 0 0 0 211 199 0 0 3
2480 2593
2526 2593
2526 2559
1 7 253 0 0 0 0 198 211 0 0 3
2513 2558
2513 2581
2480 2581
8 1 254 0 0 0 0 211 197 0 0 3
2480 2569
2500 2569
2500 2558
0 1 222 0 0 0 0 0 214 506 0 3
2199 2457
2199 2635
2247 2635
0 1 223 0 0 0 0 0 215 507 0 3
2206 2423
2206 2601
2246 2601
1 0 224 0 0 0 0 213 0 0 508 3
2246 2568
2214 2568
2214 2390
1 0 225 0 0 0 0 212 0 0 509 3
2245 2534
2221 2534
2221 2356
5 0 256 0 0 8320 0 254 0 0 489 4
2735 1922
2597 1922
2597 2409
2535 2409
0 5 257 0 0 8320 0 0 250 490 0 4
2524 2397
2605 2397
2605 2042
2734 2042
0 5 258 0 0 8320 0 0 246 491 0 4
2512 2384
2590 2384
2590 2167
2733 2167
0 5 259 0 0 12416 0 0 242 492 0 4
2497 2373
2568 2373
2568 2289
2732 2289
5 1 256 0 0 0 0 222 201 0 0 3
2478 2409
2538 2409
2538 2363
6 1 257 0 0 0 0 222 202 0 0 3
2478 2397
2525 2397
2525 2363
1 7 258 0 0 0 0 203 222 0 0 3
2512 2362
2512 2385
2478 2385
8 1 259 0 0 0 0 222 204 0 0 3
2478 2373
2499 2373
2499 2362
4 0 260 0 0 4096 0 302 0 0 495 2
1860 2268
1860 2518
5 0 260 0 0 0 0 303 0 0 495 2
1520 2263
1520 2480
0 1 260 0 0 8320 0 0 216 790 0 5
534 1769
534 2480
1824 2480
1824 2518
2418 2518
3 1 261 0 0 4224 0 208 205 0 0 4
2295 2822
2386 2822
2386 2783
2435 2783
2 3 262 0 0 12416 0 205 209 0 0 4
2435 2771
2369 2771
2369 2788
2294 2788
3 3 263 0 0 4224 0 207 205 0 0 4
2293 2755
2386 2755
2386 2759
2435 2759
4 3 264 0 0 12416 0 205 206 0 0 4
2435 2747
2405 2747
2405 2721
2293 2721
2 9 265 0 0 8320 0 210 205 0 0 3
2457 2696
2459 2696
2459 2711
3 1 266 0 0 4224 0 214 211 0 0 4
2292 2644
2383 2644
2383 2605
2432 2605
2 3 267 0 0 12416 0 211 215 0 0 4
2432 2593
2366 2593
2366 2610
2291 2610
3 3 268 0 0 4224 0 213 211 0 0 4
2291 2577
2383 2577
2383 2581
2432 2581
4 3 269 0 0 12416 0 211 212 0 0 4
2432 2569
2402 2569
2402 2543
2290 2543
2 9 270 0 0 8320 0 216 211 0 0 3
2454 2518
2456 2518
2456 2533
0 2 222 0 0 0 0 0 225 603 0 5
1944 2425
1944 2477
2037 2477
2037 2457
2245 2457
2 0 223 0 0 4096 0 226 0 0 636 2
2244 2423
1991 2423
2 0 224 0 0 4096 0 224 0 0 604 2
2244 2390
1998 2390
2 0 225 0 0 4096 0 223 0 0 635 2
2243 2356
2004 2356
0 1 16 0 0 0 0 0 225 639 0 3
1959 2399
1959 2439
2245 2439
1 0 15 0 0 0 0 226 0 0 605 2
2244 2405
1965 2405
1 0 14 0 0 0 0 224 0 0 638 2
2244 2372
1971 2372
1 0 13 0 0 0 0 223 0 0 637 2
2243 2338
1978 2338
3 1 271 0 0 4224 0 225 222 0 0 4
2290 2448
2381 2448
2381 2409
2430 2409
2 3 272 0 0 12416 0 222 226 0 0 4
2430 2397
2364 2397
2364 2414
2289 2414
3 3 273 0 0 4224 0 224 222 0 0 4
2289 2381
2381 2381
2381 2385
2430 2385
4 3 274 0 0 12416 0 222 223 0 0 4
2430 2373
2400 2373
2400 2347
2288 2347
4 0 275 0 0 4096 0 303 0 0 520 2
1511 2263
1511 2451
4 0 275 0 0 0 0 304 0 0 520 2
1170 2259
1170 2419
0 1 275 0 0 8320 0 0 221 791 0 13
540 1778
540 2419
1200 2419
1200 2451
1542 2451
1542 2475
1831 2475
1831 2487
1878 2487
1878 2472
2025 2472
2025 2325
2418 2325
2 9 276 0 0 4224 0 221 222 0 0 2
2454 2325
2454 2337
9 3 277 0 0 8320 0 262 227 0 0 4
2884 2107
2884 2164
2961 2164
2961 2228
0 4 278 0 0 4224 0 0 251 616 0 3
2396 2199
2514 2199
2514 2195
3 0 279 0 0 4224 0 251 0 0 615 2
2514 2207
2405 2207
0 2 280 0 0 12288 0 0 251 614 0 4
2421 2216
2458 2216
2458 2219
2514 2219
1 0 281 0 0 4096 0 251 0 0 613 3
2514 2231
2433 2231
2433 2225
0 4 282 0 0 4224 0 0 252 621 0 4
2395 2033
2491 2033
2491 2038
2515 2038
3 0 283 0 0 12288 0 252 0 0 620 5
2515 2050
2464 2050
2464 2045
2393 2045
2393 2041
0 2 284 0 0 8192 0 0 252 619 0 3
2413 2050
2413 2062
2515 2062
0 1 285 0 0 8192 0 0 252 618 0 3
2424 2059
2424 2074
2515 2074
5 6 286 0 0 8320 0 251 254 0 0 4
2562 2231
2580 2231
2580 1913
2735 1913
6 6 287 0 0 8320 0 250 251 0 0 4
2734 2033
2585 2033
2585 2219
2562 2219
7 6 288 0 0 12416 0 251 246 0 0 4
2562 2207
2573 2207
2573 2158
2733 2158
8 6 289 0 0 12416 0 251 242 0 0 4
2562 2195
2577 2195
2577 2280
2732 2280
8 7 290 0 0 8320 0 252 242 0 0 4
2563 2038
2569 2038
2569 2271
2732 2271
7 7 291 0 0 12416 0 252 246 0 0 4
2563 2050
2601 2050
2601 2149
2733 2149
6 7 292 0 0 12416 0 252 250 0 0 4
2563 2062
2583 2062
2583 2024
2734 2024
7 5 293 0 0 8320 0 254 252 0 0 4
2735 1904
2578 1904
2578 2074
2563 2074
1 0 294 0 0 4096 0 231 0 0 573 4
2559 2160
2544 2160
2544 2148
2538 2148
2 2 295 0 0 4224 0 231 234 0 0 2
2559 2124
2559 2128
0 1 296 0 0 4224 0 0 232 574 0 3
2539 1997
2554 1997
2554 1988
2 2 297 0 0 4224 0 232 235 0 0 2
2554 1952
2554 1957
3 3 298 0 0 4224 0 234 237 0 0 5
2574 2117
2574 1830
2600 1830
2600 1821
2620 1821
3 2 299 0 0 4224 0 235 237 0 0 5
2569 1946
2569 1834
2596 1834
2596 1812
2621 1812
1 0 300 0 0 4224 0 234 0 0 612 3
2544 2117
2339 2117
2339 2187
0 1 301 0 0 8320 0 0 235 617 0 3
2344 2021
2344 1946
2539 1946
1 0 302 0 0 4224 0 236 0 0 622 3
2574 1787
2336 1787
2336 1862
1 0 303 0 0 4224 0 233 0 0 575 2
2552 1821
2540 1821
2 2 304 0 0 4224 0 233 236 0 0 3
2588 1821
2588 1798
2589 1798
1 3 305 0 0 4224 0 237 236 0 0 3
2620 1803
2620 1787
2604 1787
1 4 306 0 0 8320 0 238 237 0 0 4
2921 2020
2871 2020
2871 1812
2666 1812
8 8 307 0 0 8320 0 253 242 0 0 4
2564 1863
2594 1863
2594 2262
2732 2262
7 8 308 0 0 8320 0 253 246 0 0 4
2564 1875
2588 1875
2588 2140
2733 2140
6 8 309 0 0 12416 0 253 250 0 0 4
2564 1887
2583 1887
2583 2015
2734 2015
8 5 310 0 0 4224 0 254 253 0 0 4
2735 1895
2579 1895
2579 1899
2564 1899
0 4 311 0 0 4096 0 0 253 626 0 4
2396 1871
2489 1871
2489 1863
2516 1863
3 0 312 0 0 4096 0 253 0 0 625 4
2516 1875
2414 1875
2414 1880
2409 1880
2 0 313 0 0 8192 0 253 0 0 624 3
2516 1887
2516 1889
2419 1889
1 0 314 0 0 8192 0 253 0 0 623 3
2516 1899
2516 1898
2434 1898
4 3 315 0 0 8320 0 262 239 0 0 4
2860 2077
2856 2077
2856 2352
2854 2352
3 3 316 0 0 8320 0 262 243 0 0 4
2860 2065
2848 2065
2848 2226
2847 2226
3 2 317 0 0 4224 0 247 262 0 0 3
2843 2102
2843 2053
2860 2053
2 3 318 0 0 4224 0 239 240 0 0 3
2808 2361
2780 2361
2780 2352
1 2 319 0 0 4224 0 239 241 0 0 2
2808 2343
2808 2330
1 9 320 0 0 4224 0 241 242 0 0 2
2808 2294
2788 2294
2 3 321 0 0 4224 0 243 244 0 0 3
2801 2235
2780 2235
2780 2229
1 2 322 0 0 4224 0 243 245 0 0 4
2801 2217
2801 2212
2799 2212
2799 2208
1 9 323 0 0 4224 0 245 246 0 0 2
2799 2172
2789 2172
2 3 324 0 0 4224 0 247 248 0 0 3
2797 2111
2781 2111
2781 2107
1 2 325 0 0 4224 0 247 249 0 0 4
2797 2093
2797 2089
2793 2089
2793 2086
1 9 326 0 0 4224 0 249 250 0 0 3
2793 2050
2790 2050
2790 2047
3 1 327 0 0 8320 0 257 262 0 0 3
2850 1976
2860 1976
2860 2041
9 3 294 0 0 4224 0 251 263 0 0 2
2538 2159
2538 2138
9 3 296 0 0 0 0 252 264 0 0 4
2539 2002
2539 1995
2543 1995
2543 1989
9 3 303 0 0 0 0 253 265 0 0 4
2540 1827
2540 1818
2546 1818
2546 1810
0 2 328 0 0 4096 0 0 263 588 0 3
2449 1800
2449 2147
2487 2147
0 1 329 0 0 4096 0 0 263 579 0 3
2471 2109
2471 2129
2487 2129
1 0 330 0 0 8192 0 264 0 0 587 3
2492 1980
2486 1980
2486 1966
3 2 329 0 0 4224 0 228 264 0 0 4
2086 2109
2484 2109
2484 1998
2492 1998
2 3 331 0 0 4224 0 257 256 0 0 3
2804 1985
2783 1985
2783 1981
1 2 332 0 0 4224 0 257 255 0 0 3
2804 1967
2799 1967
2799 1966
1 9 333 0 0 8320 0 255 254 0 0 3
2799 1930
2799 1927
2791 1927
8 1 334 0 0 8320 0 262 261 0 0 3
2908 2077
2954 2077
2954 2020
7 1 335 0 0 4224 0 262 260 0 0 3
2908 2065
2967 2065
2967 2020
6 1 336 0 0 4224 0 262 259 0 0 3
2908 2053
2980 2053
2980 2020
5 1 337 0 0 4224 0 262 258 0 0 3
2908 2041
2993 2041
2993 2020
3 2 330 0 0 4224 0 229 265 0 0 3
2088 1966
2495 1966
2495 1819
3 1 328 0 0 4224 0 230 265 0 0 4
2087 1800
2449 1800
2449 1801
2495 1801
8 0 218 0 0 0 0 266 0 0 597 3
2240 2243
2150 2243
2150 2194
0 7 219 0 0 0 0 0 266 634 0 3
2155 2182
2155 2234
2240 2234
0 6 220 0 0 0 0 0 266 598 0 3
2160 2170
2160 2225
2240 2225
0 5 221 0 0 0 0 0 266 633 0 3
2164 2158
2164 2216
2240 2216
4 0 16 0 0 0 0 266 0 0 639 3
2240 2207
2210 2207
2210 1880
3 0 15 0 0 0 0 266 0 0 605 3
2240 2198
2215 2198
2215 1871
2 0 14 0 0 0 0 266 0 0 638 3
2240 2189
2222 2189
2222 1865
1 0 13 0 0 0 0 266 0 0 637 3
2240 2180
2227 2180
2227 1853
8 0 218 0 0 0 0 272 0 0 736 5
2240 2077
2201 2077
2201 2194
1894 2194
1894 2044
6 0 220 0 0 0 0 272 0 0 734 5
2240 2059
2180 2059
2180 2170
1907 2170
1907 2068
0 8 222 0 0 0 0 0 283 603 0 3
2165 2041
2165 1916
2239 1916
0 7 223 0 0 0 0 0 283 636 0 3
2153 2032
2153 1907
2239 1907
0 6 224 0 0 0 0 0 283 604 0 3
2140 2026
2140 1898
2239 1898
5 0 225 0 0 0 0 283 0 0 635 3
2239 1889
2132 1889
2132 2014
0 4 222 0 0 8320 0 0 272 695 0 7
1562 2013
1562 2425
1984 2425
1984 2050
2154 2050
2154 2041
2240 2041
0 2 224 0 0 8320 0 0 272 693 0 6
1574 2097
1574 2437
1998 2437
1998 2026
2240 2026
2240 2023
3 0 15 0 0 0 0 283 0 0 698 7
2239 1871
2115 1871
2115 1877
1965 1877
1965 2406
1226 2406
1226 2061
2 0 338 0 0 4096 0 228 0 0 607 2
2040 2118
2020 2118
0 2 338 0 0 20608 0 0 230 627 0 7
1835 2456
1835 2478
1871 2478
1871 2466
2020 2466
2020 1809
2041 1809
1 0 339 0 0 4096 0 228 0 0 609 2
2040 2100
2014 2100
0 2 339 0 0 20480 0 0 229 629 0 7
1841 2449
1841 2472
1863 2472
1863 2457
2014 2457
2014 1975
2042 1975
1 0 340 0 0 4096 0 229 0 0 611 2
2042 1957
2009 1957
0 1 340 0 0 32896 0 0 230 631 0 10
1218 2417
1224 2417
1224 2444
1551 2444
1551 2465
1857 2465
1857 2450
2009 2450
2009 1791
2041 1791
14 1 300 0 0 0 0 266 267 0 0 4
2304 2180
2323 2180
2323 2187
2360 2187
10 1 281 0 0 4224 0 266 268 0 0 3
2304 2225
2436 2225
2436 2188
11 1 280 0 0 4224 0 266 269 0 0 3
2304 2216
2423 2216
2423 2188
12 1 279 0 0 0 0 266 270 0 0 3
2304 2207
2410 2207
2410 2187
13 1 278 0 0 0 0 266 271 0 0 5
2304 2198
2303 2198
2303 2199
2397 2199
2397 2187
14 1 301 0 0 0 0 272 273 0 0 4
2304 2014
2323 2014
2323 2021
2360 2021
10 1 285 0 0 4224 0 272 274 0 0 3
2304 2059
2436 2059
2436 2021
11 1 284 0 0 4224 0 272 275 0 0 3
2304 2050
2423 2050
2423 2022
12 1 283 0 0 4224 0 272 276 0 0 3
2304 2041
2410 2041
2410 2022
13 1 282 0 0 0 0 272 277 0 0 5
2304 2032
2303 2032
2303 2033
2397 2033
2397 2022
14 1 302 0 0 0 0 283 282 0 0 4
2303 1853
2322 1853
2322 1862
2359 1862
10 1 314 0 0 4224 0 283 281 0 0 3
2303 1898
2435 1898
2435 1864
11 1 313 0 0 4224 0 283 280 0 0 3
2303 1889
2422 1889
2422 1864
12 1 312 0 0 4224 0 283 279 0 0 3
2303 1880
2409 1880
2409 1864
13 1 311 0 0 12416 0 283 278 0 0 5
2303 1871
2302 1871
2302 1871
2396 1871
2396 1864
0 3 338 0 0 0 0 0 302 628 0 7
1158 2413
1206 2413
1206 2436
1556 2436
1556 2456
1851 2456
1851 2268
0 3 338 0 0 0 0 0 304 792 0 4
544 1787
544 2413
1161 2413
1161 2259
0 2 339 0 0 0 0 0 302 630 0 5
1502 2429
1562 2429
1562 2449
1842 2449
1842 2268
0 3 339 0 0 8320 0 0 303 793 0 6
550 1796
550 2407
1213 2407
1213 2429
1502 2429
1502 2263
0 2 340 0 0 0 0 0 303 632 0 5
1150 2401
1218 2401
1218 2424
1493 2424
1493 2263
0 2 340 0 0 0 0 0 304 794 0 4
556 1805
556 2401
1152 2401
1152 2259
5 0 221 0 0 0 0 272 0 0 733 5
2240 2050
2170 2050
2170 2158
1915 2158
1915 2080
0 7 219 0 0 0 0 0 272 735 0 5
1900 2056
1900 2182
2190 2182
2190 2068
2240 2068
0 1 225 0 0 12416 0 0 272 692 0 5
1580 2137
1580 2443
2004 2443
2004 2014
2240 2014
0 3 223 0 0 8320 0 0 272 694 0 7
1568 2058
1568 2431
1991 2431
1991 2038
2120 2038
2120 2032
2240 2032
0 1 13 0 0 0 0 0 283 696 0 5
1237 2153
1237 2420
1978 2420
1978 1853
2239 1853
0 2 14 0 0 0 0 0 283 697 0 6
1231 2105
1231 2413
1971 2413
1971 1865
2239 1865
2239 1862
0 4 16 0 0 0 0 0 283 699 0 7
1222 2022
1222 2399
1959 2399
1959 1889
2124 1889
2124 1880
2239 1880
2 0 341 0 0 4096 0 306 0 0 641 2
1034 2332
1034 2391
0 1 341 0 0 8320 0 0 302 795 0 4
564 1814
564 2391
1833 2391
1833 2268
1 0 342 0 0 4096 0 313 0 0 683 2
1097 2176
1097 2190
1 0 343 0 0 8192 0 284 0 0 752 3
1147 1555
1177 1555
1177 1677
0 2 344 0 0 8320 0 0 284 645 0 5
835 1575
835 1529
1073 1529
1073 1555
1111 1555
2 1 344 0 0 0 0 286 285 0 0 4
850 1575
835 1575
835 1595
848 1595
1 1 345 0 0 4224 0 10 286 0 0 2
792 1557
850 1557
1 2 346 0 0 4224 0 9 285 0 0 2
794 1613
848 1613
0 1 347 0 0 4096 0 0 303 649 0 2
1484 2380
1484 2263
2 0 347 0 0 8320 0 308 0 0 796 4
1725 2343
1725 2380
573 2380
573 1828
0 1 348 0 0 4224 0 0 290 700 0 4
1814 2080
1814 2039
1802 2039
1802 2030
0 1 349 0 0 4096 0 0 289 701 0 4
1822 2068
1822 2034
1815 2034
1815 2030
0 1 350 0 0 8192 0 0 288 702 0 3
1829 2056
1828 2056
1828 2030
0 1 351 0 0 4096 0 0 287 703 0 4
1836 2044
1836 2036
1841 2036
1841 2030
0 1 352 0 0 4224 0 0 291 704 0 5
1479 2082
1479 2041
1471 2041
1471 2029
1465 2029
0 1 353 0 0 4224 0 0 292 705 0 4
1488 2070
1488 2036
1478 2036
1478 2029
0 1 354 0 0 4096 0 0 293 706 0 3
1495 2058
1495 2029
1491 2029
0 1 355 0 0 4096 0 0 294 707 0 4
1500 2046
1500 2034
1504 2034
1504 2029
0 1 356 0 0 4224 0 0 298 708 0 4
1130 2085
1130 2038
1118 2038
1118 2028
0 1 357 0 0 4224 0 0 297 709 0 4
1136 2073
1136 2032
1131 2032
1131 2028
0 1 358 0 0 4096 0 0 296 710 0 4
1140 2061
1140 2034
1144 2034
1144 2028
0 1 359 0 0 8192 0 0 295 711 0 4
1143 2049
1143 2038
1157 2038
1157 2028
1 0 360 0 0 4096 0 304 0 0 663 4
1143 2259
1143 2351
1144 2351
1144 2371
2 0 360 0 0 8320 0 310 0 0 797 4
1383 2333
1383 2371
582 2371
582 1845
2 1 361 0 0 8320 0 299 308 0 0 5
1550 1859
1947 1859
1947 2356
1716 2356
1716 2343
2 1 362 0 0 12416 0 300 310 0 0 6
1263 1844
1263 1843
909 1843
909 2364
1374 2364
1374 2333
1 2 363 0 0 12416 0 306 301 0 0 4
1025 2332
1025 2354
901 2354
901 1827
0 1 364 0 0 8192 0 0 299 716 0 3
1565 1802
1550 1802
1550 1823
0 1 365 0 0 4224 0 0 301 718 0 2
1026 1791
901 1791
1 0 366 0 0 4096 0 300 0 0 717 2
1263 1808
1263 1810
9 9 367 0 0 4224 0 302 314 0 0 2
1864 2212
1864 2116
9 9 368 0 0 4224 0 303 315 0 0 4
1515 2207
1515 2133
1528 2133
1528 2118
9 9 369 0 0 4224 0 304 316 0 0 2
1174 2203
1174 2121
2 2 370 0 0 4224 0 307 311 0 0 3
1747 2246
1747 2164
1771 2164
2 2 371 0 0 4224 0 309 312 0 0 3
1405 2236
1405 2151
1436 2151
2 2 372 0 0 4224 0 305 313 0 0 3
1056 2235
1056 2161
1086 2161
1 9 373 0 0 4224 0 305 306 0 0 2
1056 2271
1056 2276
1 9 374 0 0 4224 0 307 308 0 0 2
1747 2282
1747 2287
1 9 375 0 0 4224 0 309 310 0 0 2
1405 2272
1405 2277
1 0 342 0 0 4096 0 312 0 0 683 2
1447 2166
1447 2190
3 9 376 0 0 4224 0 311 330 0 0 3
1782 2149
1782 2110
1781 2110
9 3 377 0 0 4224 0 329 312 0 0 2
1447 2112
1447 2136
3 9 378 0 0 4224 0 313 328 0 0 2
1097 2146
1097 2115
1 3 342 0 0 8320 0 311 346 0 0 3
1782 2179
1782 2190
662 2190
8 1 379 0 0 4224 0 343 338 0 0 3
1601 1835
1601 2119
1669 2119
7 1 380 0 0 4224 0 343 337 0 0 3
1613 1835
1613 2079
1670 2079
6 1 381 0 0 4224 0 343 336 0 0 3
1625 1835
1625 2040
1671 2040
1 5 382 0 0 8320 0 335 343 0 0 3
1672 1995
1637 1995
1637 1835
8 1 383 0 0 12416 0 344 334 0 0 5
1335 1834
1335 1888
1274 1888
1274 2135
1320 2135
7 1 384 0 0 12416 0 344 333 0 0 5
1347 1834
1347 1897
1287 1897
1287 2087
1320 2087
6 1 385 0 0 12416 0 344 332 0 0 5
1359 1834
1359 1907
1301 1907
1301 2040
1321 2040
5 1 386 0 0 4224 0 344 331 0 0 5
1371 1834
1371 1916
1311 1916
1311 1993
1320 1993
8 2 225 0 0 0 0 315 338 0 0 4
1552 2082
1557 2082
1557 2137
1669 2137
7 2 224 0 0 0 0 315 337 0 0 4
1552 2070
1565 2070
1565 2097
1670 2097
6 2 223 0 0 0 0 315 336 0 0 2
1552 2058
1671 2058
5 2 222 0 0 0 0 315 335 0 0 4
1552 2046
1555 2046
1555 2013
1672 2013
8 2 13 0 0 0 0 316 334 0 0 3
1198 2085
1198 2153
1320 2153
7 2 14 0 0 0 0 316 333 0 0 4
1198 2073
1209 2073
1209 2105
1320 2105
2 6 15 0 0 0 0 332 316 0 0 3
1321 2058
1321 2061
1198 2061
5 2 16 0 0 0 0 316 331 0 0 5
1198 2049
1204 2049
1204 2022
1320 2022
1320 2011
4 8 348 0 0 0 0 314 330 0 0 2
1840 2080
1805 2080
3 7 349 0 0 4224 0 314 330 0 0 2
1840 2068
1805 2068
2 6 350 0 0 4224 0 314 330 0 0 2
1840 2056
1805 2056
1 5 351 0 0 4224 0 314 330 0 0 2
1840 2044
1805 2044
4 8 352 0 0 0 0 315 329 0 0 2
1504 2082
1471 2082
3 7 353 0 0 0 0 315 329 0 0 2
1504 2070
1471 2070
2 6 354 0 0 4224 0 315 329 0 0 2
1504 2058
1471 2058
1 5 355 0 0 4224 0 315 329 0 0 2
1504 2046
1471 2046
4 8 356 0 0 0 0 316 328 0 0 2
1150 2085
1121 2085
3 7 357 0 0 0 0 316 328 0 0 2
1150 2073
1121 2073
2 6 358 0 0 4224 0 316 328 0 0 2
1150 2061
1121 2061
1 5 359 0 0 4224 0 316 328 0 0 2
1150 2049
1121 2049
1 0 387 0 0 4096 0 317 0 0 729 2
1527 1626
1528 1626
1 0 388 0 0 0 0 318 0 0 730 2
1440 1628
1440 1628
1 0 389 0 0 4096 0 319 0 0 731 2
1356 1625
1357 1625
1 0 390 0 0 4096 0 320 0 0 732 2
1259 1627
1260 1627
3 9 364 0 0 12416 0 327 343 0 0 5
1041 1659
1073 1659
1073 1752
1565 1752
1565 1811
3 9 366 0 0 12416 0 326 344 0 0 6
1040 1617
1066 1617
1066 1758
1244 1758
1244 1810
1299 1810
9 3 365 0 0 0 0 345 325 0 0 5
1026 1808
1026 1696
1060 1696
1060 1577
1041 1577
1 0 391 0 0 4096 0 322 0 0 721 3
949 1586
928 1586
928 1605
2 0 391 0 0 4096 0 326 0 0 721 2
989 1626
928 1626
1 3 391 0 0 8320 0 324 285 0 0 4
949 1668
928 1668
928 1604
894 1604
1 0 392 0 0 4096 0 323 0 0 724 2
951 1608
936 1608
1 0 392 0 0 8192 0 321 0 0 724 3
949 1568
949 1567
929 1567
1 3 392 0 0 8320 0 327 286 0 0 6
990 1650
936 1650
936 1567
929 1567
929 1566
896 1566
1 2 393 0 0 4224 0 326 323 0 0 2
989 1608
987 1608
2 2 394 0 0 4224 0 325 322 0 0 2
990 1586
985 1586
1 2 395 0 0 4224 0 325 321 0 0 2
990 1568
985 1568
2 2 396 0 0 4224 0 324 327 0 0 2
985 1668
990 1668
3 0 387 0 0 4096 0 342 0 0 758 2
1528 1622
1528 1778
3 0 388 0 0 4096 0 341 0 0 760 2
1440 1615
1440 1772
3 0 389 0 0 4096 0 340 0 0 762 2
1357 1616
1357 1767
3 0 390 0 0 4096 0 339 0 0 764 2
1260 1619
1260 1763
3 8 221 0 0 8320 0 75 314 0 0 5
922 1971
922 1929
1941 1929
1941 2080
1888 2080
3 7 220 0 0 8320 0 74 314 0 0 5
962 1973
962 1936
1934 1936
1934 2068
1888 2068
3 6 219 0 0 8320 0 73 314 0 0 5
998 1972
998 1946
1927 1946
1927 2056
1888 2056
3 5 218 0 0 8320 0 72 314 0 0 5
1035 1970
1035 1955
1922 1955
1922 2044
1888 2044
4 4 397 0 0 8320 0 75 328 0 0 3
931 2017
931 2085
1073 2085
4 3 398 0 0 8320 0 74 328 0 0 3
971 2019
971 2073
1073 2073
2 4 399 0 0 4224 0 328 73 0 0 3
1073 2061
1007 2061
1007 2018
1 4 400 0 0 8320 0 328 72 0 0 3
1073 2049
1044 2049
1044 2016
4 3 401 0 0 4224 0 330 338 0 0 3
1757 2080
1757 2128
1715 2128
3 3 402 0 0 12416 0 330 337 0 0 4
1757 2068
1740 2068
1740 2088
1716 2088
2 3 403 0 0 12416 0 330 336 0 0 4
1757 2056
1747 2056
1747 2049
1717 2049
3 1 404 0 0 8320 0 335 330 0 0 3
1718 2004
1757 2004
1757 2044
4 3 405 0 0 8320 0 329 334 0 0 4
1423 2082
1415 2082
1415 2144
1366 2144
3 3 406 0 0 4224 0 329 333 0 0 4
1423 2070
1392 2070
1392 2096
1366 2096
2 3 407 0 0 4224 0 329 332 0 0 4
1423 2058
1391 2058
1391 2049
1367 2049
1 3 408 0 0 8320 0 329 331 0 0 3
1423 2046
1423 2002
1366 2002
2 0 343 0 0 0 0 341 0 0 752 2
1429 1600
1429 1677
2 0 343 0 0 0 0 340 0 0 752 2
1346 1601
1346 1677
2 0 343 0 0 0 0 339 0 0 752 2
1249 1604
1249 1677
2 1 343 0 0 8320 0 342 11 0 0 3
1517 1607
1517 1677
1171 1677
1 1 409 0 0 4224 0 15 342 0 0 2
1528 1585
1528 1592
1 1 410 0 0 4224 0 14 341 0 0 2
1440 1578
1440 1585
1 1 411 0 0 4224 0 13 340 0 0 2
1357 1579
1357 1586
1 1 412 0 0 4224 0 12 339 0 0 2
1260 1582
1260 1589
1 0 387 0 0 0 0 344 0 0 758 2
1371 1786
1371 1778
1 1 387 0 0 8320 0 345 343 0 0 4
1098 1784
1098 1778
1637 1778
1637 1787
2 0 388 0 0 0 0 344 0 0 760 2
1359 1786
1359 1772
2 2 388 0 0 8320 0 345 343 0 0 4
1086 1784
1086 1772
1625 1772
1625 1787
3 0 389 0 0 0 0 344 0 0 762 2
1347 1786
1347 1767
3 3 389 0 0 8320 0 343 345 0 0 4
1613 1787
1613 1767
1074 1767
1074 1784
4 0 390 0 0 0 0 344 0 0 764 2
1335 1786
1335 1763
4 4 390 0 0 8320 0 345 343 0 0 4
1062 1784
1062 1763
1601 1763
1601 1787
3 0 123 0 0 0 0 350 0 0 1102 2
746 1023
746 1092
3 0 124 0 0 0 0 349 0 0 1103 2
783 1023
783 1080
3 0 125 0 0 0 0 347 0 0 1104 2
822 1023
822 1068
3 0 126 0 0 0 0 348 0 0 1105 2
859 1023
859 1056
0 2 92 0 0 0 0 0 348 770 0 3
811 1033
848 1033
848 1008
2 0 92 0 0 0 0 347 0 0 771 3
811 1008
811 1034
770 1034
0 2 92 0 0 0 0 0 349 772 0 4
721 1008
721 1034
772 1034
772 1008
0 2 92 0 0 0 0 0 350 1106 0 3
640 1148
640 1008
735 1008
1 1 413 0 0 4224 0 348 17 0 0 2
859 993
859 982
1 1 414 0 0 4224 0 347 16 0 0 2
822 993
822 982
1 1 415 0 0 4224 0 349 18 0 0 2
783 993
783 982
1 1 416 0 0 4224 0 350 19 0 0 2
746 993
746 982
4 0 417 0 0 8320 0 365 0 0 798 4
385 1742
369 1742
369 1485
538 1485
0 3 418 0 0 8320 0 0 365 799 0 4
519 1473
373 1473
373 1733
385 1733
2 0 419 0 0 8320 0 365 0 0 800 4
385 1724
379 1724
379 1461
499 1461
0 1 420 0 0 8320 0 0 365 801 0 3
480 1449
385 1449
385 1715
1 5 421 0 0 4224 0 20 365 0 0 4
329 1748
371 1748
371 1769
385 1769
22 1 71 0 0 0 0 365 353 0 0 4
449 1697
564 1697
564 1604
586 1604
21 1 78 0 0 0 0 365 354 0 0 4
449 1706
555 1706
555 1620
587 1620
20 1 102 0 0 0 0 365 352 0 0 4
449 1715
575 1715
575 1636
587 1636
19 1 198 0 0 0 0 365 351 0 0 4
449 1724
570 1724
570 1652
587 1652
18 1 200 0 0 0 0 365 357 0 0 4
449 1733
559 1733
559 1669
586 1669
17 1 201 0 0 0 0 365 358 0 0 4
449 1742
580 1742
580 1685
587 1685
16 1 226 0 0 0 0 365 356 0 0 4
449 1751
565 1751
565 1701
587 1701
15 1 255 0 0 0 0 365 355 0 0 4
449 1760
575 1760
575 1717
587 1717
14 1 260 0 0 0 0 365 360 0 0 4
449 1769
570 1769
570 1733
587 1733
13 1 275 0 0 0 0 365 359 0 0 4
449 1778
580 1778
580 1748
587 1748
12 1 338 0 0 0 0 365 361 0 0 4
449 1787
575 1787
575 1764
587 1764
11 1 339 0 0 0 0 365 362 0 0 4
449 1796
580 1796
580 1780
587 1780
10 1 340 0 0 0 0 365 363 0 0 4
449 1805
580 1805
580 1798
587 1798
1 9 341 0 0 0 0 367 365 0 0 2
587 1814
449 1814
1 8 347 0 0 0 0 366 365 0 0 4
587 1828
464 1828
464 1823
449 1823
7 1 360 0 0 0 0 365 364 0 0 4
449 1832
464 1832
464 1845
587 1845
1 5 417 0 0 0 0 371 536 0 0 3
538 1439
538 1485
555 1485
6 1 418 0 0 0 0 536 370 0 0 3
555 1473
518 1473
518 1439
1 7 419 0 0 0 0 369 536 0 0 3
499 1439
499 1461
555 1461
1 8 420 0 0 0 0 368 536 0 0 3
480 1439
480 1449
555 1449
1 0 67 0 0 0 0 372 0 0 806 2
2922 1714
2922 1759
0 1 68 0 0 0 0 0 373 807 0 2
2902 1747
2902 1714
1 0 69 0 0 0 0 374 0 0 808 2
2883 1714
2883 1735
1 0 70 0 0 0 0 376 0 0 809 2
2864 1714
2864 1723
5 1 67 0 0 4224 0 375 536 0 0 4
3056 1759
1718 1759
1718 1485
603 1485
6 2 68 0 0 4224 0 375 536 0 0 4
3056 1747
1725 1747
1725 1473
603 1473
7 3 69 0 0 4224 0 375 536 0 0 4
3056 1735
1732 1735
1732 1461
603 1461
8 4 70 0 0 4224 0 375 536 0 0 4
3056 1723
1740 1723
1740 1449
603 1449
0 3 153 0 0 0 0 0 397 0 0 5
1828 1661
1828 1662
1823 1662
1823 1661
1815 1661
3 4 422 0 0 8320 0 395 375 0 0 4
3261 937
3349 937
3349 1723
3104 1723
3 3 423 0 0 8320 0 388 375 0 0 4
3272 1169
3341 1169
3341 1735
3104 1735
3 2 424 0 0 8320 0 385 375 0 0 4
3312 1393
3335 1393
3335 1747
3104 1747
1 3 425 0 0 4224 0 375 378 0 0 3
3104 1759
3310 1759
3310 1655
1 9 426 0 0 4224 0 379 381 0 0 2
3259 1578
3264 1578
1 9 427 0 0 4224 0 384 382 0 0 2
3245 1336
3247 1336
1 9 428 0 0 4224 0 377 380 0 0 2
3249 1484
3252 1484
2 1 429 0 0 8320 0 377 378 0 0 3
3285 1484
3319 1484
3319 1609
2 2 430 0 0 8320 0 379 378 0 0 3
3295 1578
3301 1578
3301 1609
8 8 431 0 0 8320 0 417 381 0 0 5
2981 1545
2981 1634
3166 1634
3166 1610
3208 1610
8 7 432 0 0 8320 0 423 381 0 0 5
2655 1549
2655 1640
3187 1640
3187 1601
3208 1601
8 6 433 0 0 8320 0 429 381 0 0 5
2367 1547
2367 1645
3184 1645
3184 1592
3208 1592
8 5 434 0 0 8320 0 435 381 0 0 5
2076 1550
2076 1652
3181 1652
3181 1583
3208 1583
7 4 435 0 0 12288 0 0 381 837 0 5
2987 1312
2987 1347
3165 1347
3165 1574
3208 1574
8 3 436 0 0 16512 0 447 381 0 0 7
2661 1314
2661 1312
2660 1312
2660 1349
3186 1349
3186 1565
3208 1565
8 2 437 0 0 8320 0 453 381 0 0 5
2373 1311
2373 1351
3171 1351
3171 1556
3208 1556
8 1 438 0 0 8320 0 459 381 0 0 5
2082 1314
2082 1360
3187 1360
3187 1547
3208 1547
8 8 439 0 0 12416 0 465 380 0 0 5
2990 1096
2990 1124
3152 1124
3152 1516
3196 1516
8 7 440 0 0 8320 0 471 380 0 0 5
2664 1099
2664 1129
3145 1129
3145 1507
3196 1507
8 6 441 0 0 8320 0 477 380 0 0 5
2376 1094
2376 1133
3135 1133
3135 1498
3196 1498
8 5 442 0 0 8320 0 483 380 0 0 5
2085 1099
2085 1137
3128 1137
3128 1489
3196 1489
8 4 443 0 0 12416 0 489 380 0 0 5
2980 872
2980 894
3136 894
3136 1480
3196 1480
8 3 444 0 0 12416 0 495 380 0 0 5
2666 878
2666 901
3126 901
3126 1471
3196 1471
8 2 445 0 0 8320 0 501 380 0 0 5
2385 874
2385 905
3129 905
3129 1462
3196 1462
8 1 446 0 0 8320 0 507 380 0 0 5
2084 880
2084 910
3120 910
3120 1453
3196 1453
4 6 447 0 0 8320 0 391 441 0 0 5
3169 1107
3156 1107
3156 1347
2963 1347
2963 1312
8 0 435 0 0 0 0 441 0 0 846 2
2987 1312
2987 1351
2 1 448 0 0 8320 0 386 385 0 0 3
3266 1251
3321 1251
3321 1347
2 2 449 0 0 4224 0 384 385 0 0 3
3281 1336
3303 1336
3303 1347
1 9 450 0 0 4224 0 386 383 0 0 2
3230 1251
3232 1251
7 8 451 0 0 12416 0 417 382 0 0 5
2969 1545
2969 1636
3154 1636
3154 1368
3191 1368
7 7 452 0 0 8320 0 423 382 0 0 5
2643 1549
2643 1642
3175 1642
3175 1359
3191 1359
7 6 453 0 0 8320 0 429 382 0 0 5
2355 1547
2355 1647
3172 1647
3172 1350
3191 1350
7 5 454 0 0 8320 0 435 382 0 0 5
2064 1550
2064 1654
3169 1654
3169 1341
3191 1341
7 4 455 0 0 8320 0 441 382 0 0 5
2975 1312
2975 1349
3153 1349
3153 1332
3191 1332
7 3 435 0 0 12416 0 447 382 0 0 6
2649 1314
2648 1314
2648 1351
3174 1351
3174 1323
3191 1323
7 2 456 0 0 8320 0 453 382 0 0 5
2361 1311
2361 1353
3159 1353
3159 1314
3191 1314
7 1 457 0 0 8320 0 459 382 0 0 5
2070 1314
2070 1362
3175 1362
3175 1305
3191 1305
7 8 458 0 0 8320 0 465 383 0 0 5
2978 1096
2978 1126
3140 1126
3140 1283
3176 1283
7 7 459 0 0 8320 0 471 383 0 0 5
2652 1099
2652 1131
3133 1131
3133 1274
3176 1274
7 6 460 0 0 8320 0 477 383 0 0 5
2364 1094
2364 1135
3123 1135
3123 1265
3176 1265
7 5 461 0 0 8320 0 483 383 0 0 5
2073 1099
2073 1139
3116 1139
3116 1256
3176 1256
7 4 462 0 0 12416 0 489 383 0 0 5
2968 872
2968 896
3124 896
3124 1247
3176 1247
7 3 463 0 0 8320 0 495 383 0 0 5
2654 878
2654 903
3114 903
3114 1238
3176 1238
7 2 464 0 0 8320 0 501 383 0 0 5
2373 874
2373 907
3117 907
3117 1229
3176 1229
7 1 465 0 0 8320 0 507 383 0 0 5
2072 880
2072 912
3108 912
3108 1220
3176 1220
2 1 466 0 0 8320 0 387 388 0 0 3
3261 1037
3281 1037
3281 1123
2 2 467 0 0 4224 0 388 389 0 0 3
3263 1123
3263 1111
3260 1111
1 9 468 0 0 4224 0 389 391 0 0 2
3224 1111
3225 1111
1 9 469 0 0 0 0 387 390 0 0 2
3225 1037
3225 1037
6 0 470 0 0 0 0 507 0 0 890 2
2060 880
2060 880
6 0 471 0 0 0 0 501 0 0 889 2
2361 874
2361 874
6 0 472 0 0 0 0 495 0 0 888 2
2642 878
2642 878
6 0 473 0 0 0 0 489 0 0 887 2
2956 872
2956 872
6 0 474 0 0 0 0 483 0 0 886 2
2061 1099
2061 1099
6 0 475 0 0 0 0 477 0 0 885 2
2352 1094
2352 1094
6 0 476 0 0 0 0 471 0 0 884 2
2640 1099
2640 1099
6 0 477 0 0 0 0 465 0 0 883 2
2966 1096
2966 1096
6 0 478 0 0 0 0 459 0 0 882 2
2058 1314
2058 1314
6 0 479 0 0 0 0 453 0 0 881 2
2349 1311
2349 1311
6 0 480 0 0 0 0 447 0 0 880 2
2637 1314
2637 1314
6 0 481 0 0 0 0 435 0 0 879 2
2052 1550
2052 1550
6 0 482 0 0 0 0 429 0 0 878 2
2343 1547
2343 1547
6 0 483 0 0 0 0 423 0 0 877 2
2631 1549
2631 1549
6 0 484 0 0 0 0 417 0 0 876 2
2957 1545
2957 1545
5 8 484 0 0 12416 0 0 391 0 0 4
2957 1541
2957 1633
3169 1633
3169 1143
5 7 483 0 0 8320 0 0 391 0 0 5
2631 1545
2631 1639
3165 1639
3165 1134
3169 1134
5 6 482 0 0 8320 0 0 391 0 0 5
2343 1543
2343 1644
3160 1644
3160 1125
3169 1125
5 5 481 0 0 8320 0 0 391 0 0 5
2052 1546
2052 1651
3157 1651
3157 1116
3169 1116
5 3 480 0 0 8320 0 0 391 0 0 5
2637 1310
2637 1355
3152 1355
3152 1098
3169 1098
5 2 479 0 0 8320 0 0 391 0 0 5
2349 1307
2349 1361
3144 1361
3144 1089
3169 1089
5 1 478 0 0 8320 0 0 391 0 0 5
2058 1310
2058 1367
3132 1367
3132 1080
3169 1080
5 8 477 0 0 8320 0 0 390 0 0 5
2966 1092
2966 1123
3128 1123
3128 1069
3169 1069
5 7 476 0 0 8320 0 0 390 0 0 5
2640 1095
2640 1128
3121 1128
3121 1060
3169 1060
5 6 475 0 0 8320 0 0 390 0 0 5
2352 1090
2352 1132
3111 1132
3111 1051
3169 1051
5 5 474 0 0 8320 0 0 390 0 0 5
2061 1095
2061 1136
3104 1136
3104 1042
3169 1042
5 4 473 0 0 8320 0 0 390 0 0 5
2956 868
2956 893
3112 893
3112 1033
3169 1033
5 3 472 0 0 8320 0 0 390 0 0 5
2642 874
2642 900
3102 900
3102 1024
3169 1024
5 2 471 0 0 8320 0 0 390 0 0 5
2361 870
2361 904
3105 904
3105 1015
3169 1015
5 1 470 0 0 8320 0 0 390 0 0 5
2060 876
2060 909
3096 909
3096 1006
3169 1006
5 8 485 0 0 12416 0 417 392 0 0 4
2945 1545
2945 1637
3160 1637
3160 915
5 7 486 0 0 12416 0 423 392 0 0 5
2619 1549
2619 1643
3153 1643
3153 906
3160 906
5 6 487 0 0 8320 0 429 392 0 0 5
2331 1547
2331 1648
3148 1648
3148 897
3160 897
5 5 488 0 0 8320 0 435 392 0 0 5
2040 1550
2040 1655
3145 1655
3145 888
3160 888
5 4 489 0 0 12416 0 441 392 0 0 5
2951 1312
2951 1354
3136 1354
3136 879
3160 879
5 3 490 0 0 8320 0 447 392 0 0 5
2625 1314
2625 1359
3140 1359
3140 870
3160 870
5 2 491 0 0 8320 0 453 392 0 0 5
2337 1311
2337 1365
3132 1365
3132 861
3160 861
5 1 492 0 0 8320 0 459 392 0 0 5
2046 1314
2046 1371
3120 1371
3120 852
3160 852
5 8 493 0 0 12416 0 465 393 0 0 5
2954 1096
2954 1127
3116 1127
3116 843
3160 843
5 7 494 0 0 8320 0 471 393 0 0 5
2628 1099
2628 1132
3109 1132
3109 834
3160 834
5 6 495 0 0 8320 0 477 393 0 0 5
2340 1094
2340 1136
3099 1136
3099 825
3160 825
5 5 496 0 0 8320 0 483 393 0 0 5
2049 1099
2049 1140
3092 1140
3092 816
3160 816
5 4 497 0 0 8320 0 489 393 0 0 5
2944 872
2944 898
3113 898
3113 807
3160 807
5 3 498 0 0 8320 0 495 393 0 0 5
2630 878
2630 906
3105 906
3105 798
3160 798
5 2 499 0 0 8320 0 501 393 0 0 5
2349 874
2349 912
3096 912
3096 789
3160 789
5 1 500 0 0 8320 0 507 393 0 0 5
2048 880
2048 917
3088 917
3088 780
3160 780
1 9 501 0 0 0 0 394 392 0 0 2
3216 883
3216 883
2 2 502 0 0 4224 0 395 394 0 0 2
3252 891
3252 883
1 9 503 0 0 4224 0 396 393 0 0 2
3221 811
3216 811
2 1 504 0 0 8320 0 396 395 0 0 3
3257 811
3270 811
3270 891
2 0 157 0 0 8320 0 138 0 0 1199 6
3078 1472
3078 1377
1870 1377
1870 1158
1436 1158
1436 1167
2 0 159 0 0 8320 0 139 0 0 1198 6
2750 1476
2750 1389
1878 1389
1878 1142
1435 1142
1435 1150
2 0 161 0 0 8320 0 140 0 0 1197 6
2462 1471
2462 1400
1888 1400
1888 1127
1446 1127
1446 1136
2 0 163 0 0 16512 0 141 0 0 1196 6
2173 1475
2173 1411
1896 1411
1896 1110
1446 1110
1446 1120
0 2 165 0 0 16512 0 0 142 1195 0 7
1444 1102
1444 1093
1902 1093
1902 1144
3083 1144
3083 1241
3082 1241
2 0 167 0 0 12416 0 143 0 0 1194 7
2759 1240
2760 1240
2760 1155
1909 1155
1909 1077
1445 1077
1445 1086
2 0 169 0 0 12416 0 144 0 0 1193 7
2473 1241
2474 1241
2474 1166
1919 1166
1919 1063
1436 1063
1436 1070
2 0 171 0 0 16512 0 145 0 0 1192 6
2183 1245
2183 1179
1928 1179
1928 1047
1437 1047
1437 1055
0 2 173 0 0 16512 0 0 146 1191 0 7
1436 1039
1436 1031
1900 1031
1900 923
3081 923
3081 1024
3071 1024
2 0 175 0 0 8320 0 147 0 0 1190 6
2755 1028
2755 935
1911 935
1911 1015
1435 1015
1435 1023
2 0 177 0 0 12416 0 148 0 0 1189 7
2471 1020
2475 1020
2475 947
1920 947
1920 1001
1436 1001
1436 1007
2 0 179 0 0 20608 0 149 0 0 1188 7
2185 1028
2186 1028
2186 962
1927 962
1927 984
1436 984
1436 991
2 0 181 0 0 12416 0 150 0 0 1187 7
3072 802
3076 802
3076 680
1891 680
1891 762
1423 762
1423 974
2 0 183 0 0 8320 0 151 0 0 1186 6
2761 803
2761 689
1897 689
1897 770
1431 770
1431 958
2 0 186 0 0 8320 0 152 0 0 1185 6
2479 803
2479 698
1905 698
1905 781
1438 781
1438 942
1 0 153 0 0 4096 0 405 0 0 932 2
2137 1450
2210 1450
1 0 153 0 0 0 0 401 0 0 932 2
2147 1215
2210 1215
1 0 153 0 0 0 0 409 0 0 932 2
2151 999
2210 999
1 0 153 0 0 0 0 404 0 0 933 2
2430 1449
2499 1449
1 0 153 0 0 0 0 400 0 0 933 2
2439 1213
2499 1213
1 0 153 0 0 0 0 408 0 0 933 2
2441 996
2499 996
1 0 153 0 0 8192 0 509 0 0 945 3
2152 783
2210 783
2210 1661
1 0 153 0 0 8192 0 412 0 0 945 3
2450 778
2499 778
2499 1661
1 0 153 0 0 0 0 403 0 0 937 2
2721 1449
2800 1449
1 0 153 0 0 0 0 399 0 0 937 2
2726 1216
2800 1216
1 0 153 0 0 0 0 407 0 0 937 2
2725 999
2800 999
1 0 153 0 0 0 0 411 0 0 945 3
2731 779
2800 779
2800 1661
1 0 153 0 0 0 0 402 0 0 945 2
3046 1447
3126 1447
1 0 153 0 0 0 0 398 0 0 945 2
3051 1215
3126 1215
3 9 505 0 0 4224 0 398 512 0 0 2
3021 1215
3017 1215
3 9 506 0 0 4224 0 399 515 0 0 2
2696 1216
2691 1216
3 9 507 0 0 4224 0 400 518 0 0 2
2409 1213
2403 1213
3 9 508 0 0 4224 0 401 521 0 0 2
2117 1215
2112 1215
1 0 153 0 0 0 0 406 0 0 945 2
3053 999
3126 999
1 0 153 0 0 12416 0 410 0 0 0 7
3040 777
3126 777
3126 1661
2206 1661
2206 1662
1858 1662
1858 1661
3 9 509 0 0 4224 0 402 513 0 0 2
3016 1447
3011 1447
3 9 510 0 0 4224 0 403 516 0 0 2
2691 1449
2685 1449
3 9 511 0 0 4224 0 404 519 0 0 2
2400 1449
2397 1449
3 9 512 0 0 4224 0 405 520 0 0 2
2107 1450
2106 1450
3 9 513 0 0 4224 0 406 511 0 0 2
3023 999
3020 999
3 9 514 0 0 4224 0 407 514 0 0 2
2695 999
2694 999
3 9 515 0 0 4224 0 408 517 0 0 2
2411 996
2406 996
3 9 516 0 0 4224 0 409 522 0 0 2
2121 999
2115 999
3 9 517 0 0 0 0 410 523 0 0 2
3010 777
3010 777
3 9 518 0 0 4224 0 411 524 0 0 2
2701 779
2696 779
3 9 519 0 0 4224 0 412 525 0 0 2
2420 778
2415 778
3 9 520 0 0 4224 0 509 533 0 0 2
2122 783
2114 783
2 9 521 0 0 4224 0 418 417 0 0 2
3014 1521
3017 1521
1 0 522 0 0 8320 0 416 0 0 963 3
2915 1480
2915 1479
2981 1479
1 0 523 0 0 8320 0 415 0 0 964 3
2901 1480
2901 1484
2969 1484
0 1 524 0 0 4224 0 0 414 965 0 3
2957 1490
2887 1490
2887 1480
1 0 525 0 0 8320 0 413 0 0 966 3
2872 1480
2872 1497
2945 1497
4 8 522 0 0 0 0 417 513 0 0 2
2981 1497
2981 1471
3 7 523 0 0 0 0 417 513 0 0 2
2969 1497
2969 1471
2 6 524 0 0 0 0 417 513 0 0 2
2957 1497
2957 1471
1 5 525 0 0 0 0 417 513 0 0 2
2945 1497
2945 1471
2 9 526 0 0 4224 0 424 423 0 0 2
2688 1525
2691 1525
1 0 527 0 0 8320 0 422 0 0 972 3
2589 1482
2589 1481
2655 1481
1 0 528 0 0 8320 0 421 0 0 973 3
2575 1482
2575 1486
2643 1486
0 1 529 0 0 4224 0 0 420 974 0 3
2631 1492
2561 1492
2561 1482
1 0 530 0 0 8320 0 419 0 0 975 3
2546 1482
2546 1499
2619 1499
4 8 527 0 0 0 0 423 516 0 0 2
2655 1501
2655 1473
3 7 528 0 0 0 0 423 516 0 0 2
2643 1501
2643 1473
2 6 529 0 0 0 0 423 516 0 0 2
2631 1501
2631 1473
1 5 530 0 0 0 0 423 516 0 0 2
2619 1501
2619 1473
2 9 531 0 0 4224 0 430 429 0 0 2
2400 1523
2403 1523
1 0 532 0 0 8320 0 428 0 0 981 3
2301 1482
2301 1481
2367 1481
1 0 533 0 0 8320 0 427 0 0 982 3
2287 1482
2287 1486
2355 1486
0 1 534 0 0 4224 0 0 426 983 0 3
2343 1492
2273 1492
2273 1482
1 0 535 0 0 8320 0 425 0 0 984 3
2258 1482
2258 1499
2331 1499
4 8 532 0 0 0 0 429 519 0 0 2
2367 1499
2367 1473
3 7 533 0 0 0 0 429 519 0 0 2
2355 1499
2355 1473
2 6 534 0 0 0 0 429 519 0 0 2
2343 1499
2343 1473
1 5 535 0 0 0 0 429 519 0 0 2
2331 1499
2331 1473
2 9 536 0 0 4224 0 436 435 0 0 2
2109 1526
2112 1526
1 0 537 0 0 8320 0 434 0 0 990 3
2010 1483
2010 1482
2076 1482
1 0 538 0 0 8320 0 433 0 0 991 3
1996 1483
1996 1487
2064 1487
0 1 539 0 0 4224 0 0 432 992 0 3
2052 1493
1982 1493
1982 1483
1 0 540 0 0 8320 0 431 0 0 993 3
1967 1483
1967 1500
2040 1500
4 8 537 0 0 0 0 435 520 0 0 2
2076 1502
2076 1474
3 7 538 0 0 0 0 435 520 0 0 2
2064 1502
2064 1474
2 6 539 0 0 0 0 435 520 0 0 2
2052 1502
2052 1474
1 5 540 0 0 0 0 435 520 0 0 2
2040 1502
2040 1474
2 9 541 0 0 4224 0 442 441 0 0 2
3020 1288
3023 1288
1 0 542 0 0 8320 0 440 0 0 999 3
2921 1248
2921 1247
2987 1247
1 0 543 0 0 8320 0 439 0 0 1000 3
2907 1248
2907 1252
2975 1252
0 1 544 0 0 4224 0 0 438 1001 0 3
2963 1258
2893 1258
2893 1248
1 0 545 0 0 8320 0 437 0 0 1002 3
2878 1248
2878 1265
2951 1265
4 8 542 0 0 0 0 441 512 0 0 2
2987 1264
2987 1239
3 7 543 0 0 0 0 441 512 0 0 2
2975 1264
2975 1239
2 6 544 0 0 0 0 441 512 0 0 2
2963 1264
2963 1239
1 5 545 0 0 0 0 441 512 0 0 4
2951 1264
2951 1265
2951 1265
2951 1239
2 9 546 0 0 4224 0 448 447 0 0 2
2694 1290
2697 1290
1 0 547 0 0 8320 0 446 0 0 1008 3
2595 1249
2595 1248
2661 1248
1 0 548 0 0 8320 0 445 0 0 1009 3
2581 1249
2581 1253
2649 1253
0 1 549 0 0 4224 0 0 444 1010 0 3
2637 1259
2567 1259
2567 1249
1 0 550 0 0 8320 0 443 0 0 1011 3
2552 1249
2552 1266
2625 1266
4 8 547 0 0 0 0 447 515 0 0 2
2661 1266
2661 1240
3 7 548 0 0 0 0 447 515 0 0 2
2649 1266
2649 1240
2 6 549 0 0 0 0 447 515 0 0 2
2637 1266
2637 1240
1 5 550 0 0 0 0 447 515 0 0 2
2625 1266
2625 1240
2 9 551 0 0 4224 0 454 453 0 0 2
2406 1287
2409 1287
1 0 552 0 0 8320 0 452 0 0 1017 3
2307 1246
2307 1245
2373 1245
1 0 553 0 0 8320 0 451 0 0 1018 3
2293 1246
2293 1250
2361 1250
0 1 554 0 0 4224 0 0 450 1019 0 3
2349 1256
2279 1256
2279 1246
1 0 555 0 0 8320 0 449 0 0 1020 3
2264 1246
2264 1263
2337 1263
4 8 552 0 0 0 0 453 518 0 0 2
2373 1263
2373 1237
3 7 553 0 0 0 0 453 518 0 0 2
2361 1263
2361 1237
2 6 554 0 0 0 0 453 518 0 0 2
2349 1263
2349 1237
1 5 555 0 0 0 0 453 518 0 0 2
2337 1263
2337 1237
2 9 556 0 0 4224 0 460 459 0 0 2
2115 1290
2118 1290
1 0 557 0 0 8320 0 458 0 0 1026 3
2016 1248
2016 1247
2082 1247
1 0 558 0 0 8320 0 457 0 0 1027 3
2002 1248
2002 1252
2070 1252
0 1 559 0 0 4224 0 0 456 1028 0 3
2058 1258
1988 1258
1988 1248
1 0 560 0 0 8320 0 455 0 0 1029 3
1973 1248
1973 1265
2046 1265
4 8 557 0 0 0 0 459 521 0 0 2
2082 1266
2082 1239
3 7 558 0 0 0 0 459 521 0 0 2
2070 1266
2070 1239
2 6 559 0 0 0 0 459 521 0 0 2
2058 1266
2058 1239
1 5 560 0 0 0 0 459 521 0 0 2
2046 1266
2046 1239
2 9 561 0 0 4224 0 466 465 0 0 2
3023 1072
3026 1072
1 0 562 0 0 8320 0 464 0 0 1035 3
2924 1032
2924 1031
2990 1031
1 0 563 0 0 8320 0 463 0 0 1036 3
2910 1032
2910 1036
2978 1036
0 1 564 0 0 4224 0 0 462 1037 0 3
2966 1042
2896 1042
2896 1032
1 0 565 0 0 8320 0 461 0 0 1038 3
2881 1032
2881 1049
2954 1049
4 8 562 0 0 0 0 465 511 0 0 2
2990 1048
2990 1023
3 7 563 0 0 0 0 465 511 0 0 2
2978 1048
2978 1023
2 6 564 0 0 0 0 465 511 0 0 2
2966 1048
2966 1023
1 5 565 0 0 0 0 465 511 0 0 4
2954 1048
2954 1049
2954 1049
2954 1023
2 9 566 0 0 4224 0 472 471 0 0 2
2697 1075
2700 1075
1 0 567 0 0 8320 0 470 0 0 1044 3
2598 1032
2598 1031
2664 1031
1 0 568 0 0 8320 0 469 0 0 1045 3
2584 1032
2584 1036
2652 1036
0 1 569 0 0 4224 0 0 468 1046 0 3
2640 1042
2570 1042
2570 1032
1 0 570 0 0 8320 0 467 0 0 1047 3
2555 1032
2555 1049
2628 1049
4 8 567 0 0 0 0 471 514 0 0 2
2664 1051
2664 1023
3 7 568 0 0 0 0 471 514 0 0 2
2652 1051
2652 1023
2 6 569 0 0 0 0 471 514 0 0 2
2640 1051
2640 1023
1 5 570 0 0 0 0 471 514 0 0 2
2628 1051
2628 1023
2 9 571 0 0 4224 0 478 477 0 0 2
2409 1070
2412 1070
1 0 572 0 0 8320 0 476 0 0 1053 3
2310 1028
2310 1027
2376 1027
1 0 573 0 0 8320 0 475 0 0 1054 3
2296 1028
2296 1032
2364 1032
0 1 574 0 0 4224 0 0 474 1055 0 3
2352 1038
2282 1038
2282 1028
1 0 575 0 0 8320 0 473 0 0 1056 3
2267 1028
2267 1045
2340 1045
4 8 572 0 0 0 0 477 517 0 0 2
2376 1046
2376 1020
3 7 573 0 0 0 0 477 517 0 0 2
2364 1046
2364 1020
2 6 574 0 0 0 0 477 517 0 0 2
2352 1046
2352 1020
1 5 575 0 0 0 0 477 517 0 0 2
2340 1046
2340 1020
2 9 576 0 0 4224 0 484 483 0 0 2
2118 1075
2121 1075
1 0 577 0 0 4224 0 482 0 0 1062 2
2019 1032
2085 1032
1 0 578 0 0 8320 0 481 0 0 1063 3
2005 1032
2005 1036
2073 1036
0 1 579 0 0 4224 0 0 480 1064 0 3
2061 1042
1991 1042
1991 1032
1 0 580 0 0 8320 0 479 0 0 1065 3
1976 1032
1976 1049
2049 1049
4 8 577 0 0 0 0 483 522 0 0 2
2085 1051
2085 1023
3 7 578 0 0 0 0 483 522 0 0 2
2073 1051
2073 1023
2 6 579 0 0 0 0 483 522 0 0 2
2061 1051
2061 1023
1 5 580 0 0 0 0 483 522 0 0 2
2049 1051
2049 1023
4 8 581 0 0 4096 0 489 523 0 0 2
2980 824
2980 801
3 7 582 0 0 4096 0 489 523 0 0 2
2968 824
2968 801
2 6 583 0 0 4096 0 489 523 0 0 2
2956 824
2956 801
1 5 584 0 0 12288 0 489 523 0 0 4
2944 824
2944 825
2944 825
2944 801
2 9 585 0 0 4224 0 490 489 0 0 2
3013 848
3016 848
1 0 581 0 0 8320 0 488 0 0 1066 3
2914 808
2914 807
2980 807
1 0 582 0 0 8320 0 487 0 0 1067 3
2900 808
2900 812
2968 812
0 1 583 0 0 4224 0 0 486 1068 0 3
2956 818
2886 818
2886 808
1 0 584 0 0 8320 0 485 0 0 1069 3
2871 808
2871 825
2944 825
2 9 586 0 0 4224 0 496 495 0 0 2
2699 854
2702 854
1 0 587 0 0 8320 0 494 0 0 1080 3
2600 811
2600 810
2666 810
1 0 588 0 0 8320 0 493 0 0 1081 3
2586 811
2586 815
2654 815
0 1 589 0 0 4224 0 0 492 1082 0 3
2642 821
2572 821
2572 811
1 0 590 0 0 8320 0 491 0 0 1083 3
2557 811
2557 828
2630 828
4 8 587 0 0 0 0 495 524 0 0 2
2666 830
2666 803
3 7 588 0 0 0 0 495 524 0 0 2
2654 830
2654 803
2 6 589 0 0 0 0 495 524 0 0 2
2642 830
2642 803
1 5 590 0 0 0 0 495 524 0 0 2
2630 830
2630 803
2 9 591 0 0 4224 0 502 501 0 0 2
2418 850
2421 850
1 0 592 0 0 8320 0 500 0 0 1089 3
2319 810
2319 809
2385 809
1 0 593 0 0 8320 0 499 0 0 1090 3
2305 810
2305 814
2373 814
0 1 594 0 0 4224 0 0 498 1091 0 3
2361 820
2291 820
2291 810
1 0 595 0 0 8320 0 497 0 0 1092 3
2276 810
2276 827
2349 827
4 8 592 0 0 0 0 501 525 0 0 2
2385 826
2385 802
3 7 593 0 0 0 0 501 525 0 0 2
2373 826
2373 802
2 6 594 0 0 0 0 501 525 0 0 2
2361 826
2361 802
1 5 595 0 0 0 0 501 525 0 0 4
2349 826
2349 827
2349 827
2349 802
4 8 596 0 0 4096 0 507 533 0 0 2
2084 832
2084 807
3 7 597 0 0 4096 0 507 533 0 0 2
2072 832
2072 807
2 6 598 0 0 4096 0 507 533 0 0 2
2060 832
2060 807
1 5 599 0 0 4096 0 507 533 0 0 2
2048 832
2048 807
2 9 600 0 0 4224 0 508 507 0 0 2
2117 856
2120 856
1 0 596 0 0 8320 0 506 0 0 1093 3
2018 814
2018 813
2084 813
1 0 597 0 0 8320 0 505 0 0 1094 3
2004 814
2004 818
2072 818
0 1 598 0 0 4224 0 0 504 1095 0 3
2060 824
1990 824
1990 814
1 0 599 0 0 8320 0 503 0 0 1096 3
1975 814
1975 831
2048 831
4 8 123 0 0 4224 0 82 510 0 0 2
935 1092
697 1092
7 3 124 0 0 4224 0 510 82 0 0 2
697 1080
935 1080
2 6 125 0 0 4224 0 82 510 0 0 2
935 1068
697 1068
5 1 126 0 0 4224 0 510 82 0 0 2
697 1056
935 1056
1 9 92 0 0 0 0 7 510 0 0 5
611 1162
640 1162
640 1148
673 1148
673 1128
4 0 601 0 0 4096 0 516 0 0 1109 2
2655 1425
2655 1384
4 0 601 0 0 0 0 519 0 0 1109 2
2367 1425
2367 1384
0 4 601 0 0 4096 0 0 520 1110 0 3
2814 1384
2076 1384
2076 1426
4 0 601 0 0 0 0 513 0 0 1179 3
2981 1423
2981 1384
2813 1384
4 0 601 0 0 0 0 515 0 0 1113 2
2661 1192
2661 1150
4 0 601 0 0 0 0 518 0 0 1113 2
2373 1189
2373 1150
0 4 601 0 0 0 0 0 521 1114 0 3
2813 1150
2082 1150
2082 1191
4 0 601 0 0 0 0 512 0 0 1179 3
2987 1191
2987 1150
2813 1150
4 0 601 0 0 0 0 514 0 0 1117 2
2664 975
2664 928
4 0 601 0 0 0 0 517 0 0 1117 2
2376 972
2376 928
0 4 601 0 0 0 0 0 522 1118 0 3
2813 928
2085 928
2085 975
4 0 601 0 0 0 0 511 0 0 1179 3
2990 975
2990 928
2813 928
4 0 601 0 0 0 0 524 0 0 1121 2
2666 755
2666 715
4 0 601 0 0 0 0 525 0 0 1121 2
2385 754
2385 715
0 4 601 0 0 0 0 0 533 1122 0 3
2814 715
2084 715
2084 759
4 0 601 0 0 0 0 523 0 0 1179 3
2980 753
2980 715
2813 715
3 0 602 0 0 4096 0 519 0 0 1124 2
2355 1425
2355 1393
0 3 602 0 0 8192 0 0 520 1126 0 4
2511 1394
2511 1393
2064 1393
2064 1426
3 0 602 0 0 0 0 516 0 0 1126 2
2643 1425
2643 1394
0 3 602 0 0 4096 0 0 513 1177 0 3
2510 1394
2969 1394
2969 1423
3 0 602 0 0 0 0 515 0 0 1128 2
2649 1192
2649 1161
0 3 602 0 0 8192 0 0 512 1130 0 4
2510 1160
2510 1161
2975 1161
2975 1191
3 0 602 0 0 0 0 518 0 0 1130 2
2361 1189
2361 1160
0 3 602 0 0 0 0 0 521 1177 0 3
2510 1160
2070 1160
2070 1191
3 0 602 0 0 0 0 514 0 0 1132 2
2652 975
2652 940
0 3 602 0 0 8192 0 0 511 1134 0 4
2510 941
2510 940
2978 940
2978 975
3 0 602 0 0 0 0 517 0 0 1134 2
2364 972
2364 941
0 3 602 0 0 0 0 0 522 1177 0 3
2510 941
2073 941
2073 975
3 0 602 0 0 0 0 524 0 0 1136 2
2654 755
2654 725
0 3 602 0 0 0 0 0 523 1138 0 4
2509 726
2509 725
2968 725
2968 753
3 0 602 0 0 0 0 525 0 0 1138 2
2373 754
2373 726
0 3 602 0 0 0 0 0 533 1177 0 3
2510 726
2072 726
2072 759
2 0 603 0 0 4096 0 516 0 0 1141 2
2631 1425
2631 1406
2 0 603 0 0 0 0 519 0 0 1141 2
2343 1425
2343 1406
0 2 603 0 0 8192 0 0 513 1142 0 4
2216 1405
2216 1406
2957 1406
2957 1423
0 2 603 0 0 0 0 0 520 1175 0 3
2217 1405
2052 1405
2052 1426
2 0 603 0 0 0 0 515 0 0 1145 2
2637 1192
2637 1173
2 0 603 0 0 0 0 518 0 0 1145 2
2349 1189
2349 1173
0 2 603 0 0 4096 0 0 512 1146 0 3
2217 1173
2963 1173
2963 1191
0 2 603 0 0 0 0 0 521 1175 0 3
2217 1173
2058 1173
2058 1191
2 0 603 0 0 0 0 514 0 0 1149 2
2640 975
2640 953
2 0 603 0 0 0 0 517 0 0 1149 2
2352 972
2352 953
0 2 603 0 0 8192 0 0 511 1150 0 4
2217 954
2217 953
2966 953
2966 975
2 0 603 0 0 0 0 522 0 0 1175 3
2061 975
2061 954
2217 954
2 0 603 0 0 0 0 524 0 0 1153 2
2642 755
2642 736
2 0 603 0 0 0 0 525 0 0 1153 2
2361 754
2361 736
0 2 603 0 0 0 0 0 523 1154 0 3
2217 736
2956 736
2956 753
0 2 603 0 0 0 0 0 533 1175 0 3
2217 736
2060 736
2060 759
1 0 604 0 0 4096 0 516 0 0 1158 2
2619 1425
2619 1418
1 0 604 0 0 0 0 519 0 0 1158 2
2331 1425
2331 1418
1 0 604 0 0 4096 0 520 0 0 1158 2
2040 1426
2040 1418
1 0 604 0 0 8192 0 513 0 0 1180 3
2945 1423
2945 1418
1933 1418
1 0 604 0 0 0 0 515 0 0 1162 2
2625 1192
2625 1184
1 0 604 0 0 0 0 518 0 0 1162 2
2337 1189
2337 1184
1 0 604 0 0 0 0 521 0 0 1162 2
2046 1191
2046 1184
1 0 604 0 0 8192 0 512 0 0 1180 3
2951 1191
2951 1184
1933 1184
1 0 604 0 0 0 0 514 0 0 1166 2
2628 975
2628 968
1 0 604 0 0 0 0 517 0 0 1166 2
2340 972
2340 968
1 0 604 0 0 0 0 522 0 0 1166 2
2049 975
2049 968
0 1 604 0 0 4224 0 0 511 1180 0 3
1933 968
2954 968
2954 975
1 0 604 0 0 0 0 533 0 0 1170 2
2048 759
2048 747
1 0 604 0 0 0 0 525 0 0 1170 2
2349 754
2349 747
1 0 604 0 0 0 0 524 0 0 1170 2
2630 755
2630 747
0 1 604 0 0 0 0 0 523 1180 0 3
1933 747
2944 747
2944 753
2 0 90 0 0 0 0 534 0 0 1174 2
1917 595
1917 628
2 0 90 0 0 0 0 526 0 0 1174 2
2202 590
2202 628
2 0 90 0 0 0 0 528 0 0 1174 2
2495 595
2495 628
0 2 90 0 0 4224 0 0 530 0 0 3
1796 628
2798 628
2798 601
3 1 603 0 0 12416 0 526 527 0 0 4
2217 579
2217 578
2217 578
2217 1584
3 1 605 0 0 4224 0 69 526 0 0 3
2174 566
2174 579
2187 579
3 1 602 0 0 12416 0 528 529 0 0 4
2510 584
2510 583
2510 583
2510 1589
3 1 606 0 0 4224 0 68 528 0 0 3
2472 567
2472 584
2480 584
3 1 601 0 0 12416 0 530 531 0 0 4
2813 590
2813 589
2813 589
2813 1595
3 1 604 0 0 0 0 534 532 0 0 3
1932 584
1933 584
1933 1590
3 1 607 0 0 8320 0 71 534 0 0 4
1962 560
1962 569
1902 569
1902 584
1 0 132 0 0 0 0 81 0 0 1183 3
959 1183
959 1301
501 1301
3 9 132 0 0 0 0 537 535 0 0 3
339 1301
527 1301
527 1122
7 1 185 0 0 0 0 538 552 0 0 3
1377 1020
1377 926
1449 926
8 1 186 0 0 0 0 538 551 0 0 4
1377 1029
1382 1029
1382 942
1450 942
9 1 183 0 0 0 0 538 553 0 0 4
1377 1038
1388 1038
1388 958
1450 958
10 1 181 0 0 0 0 538 554 0 0 4
1377 1047
1394 1047
1394 974
1450 974
11 1 179 0 0 0 0 538 548 0 0 4
1377 1056
1400 1056
1400 991
1449 991
12 1 177 0 0 0 0 538 547 0 0 4
1377 1065
1407 1065
1407 1007
1450 1007
13 1 175 0 0 0 0 538 549 0 0 4
1377 1074
1414 1074
1414 1023
1450 1023
14 1 173 0 0 0 0 538 550 0 0 4
1377 1083
1420 1083
1420 1039
1450 1039
15 1 171 0 0 0 0 538 545 0 0 4
1377 1092
1426 1092
1426 1055
1450 1055
16 1 169 0 0 0 0 538 546 0 0 4
1377 1101
1431 1101
1431 1070
1450 1070
17 1 167 0 0 0 0 538 544 0 0 4
1377 1110
1435 1110
1435 1086
1450 1086
18 1 165 0 0 0 0 538 543 0 0 4
1377 1119
1439 1119
1439 1102
1450 1102
19 1 163 0 0 0 0 538 542 0 0 4
1377 1128
1443 1128
1443 1120
1450 1120
1 20 161 0 0 0 0 539 538 0 0 4
1450 1136
1446 1136
1446 1137
1377 1137
1 21 159 0 0 0 0 540 538 0 0 3
1450 1150
1377 1150
1377 1146
22 1 157 0 0 0 0 538 541 0 0 3
1377 1155
1377 1167
1450 1167
4 8 608 0 0 4224 0 510 535 0 0 2
649 1092
551 1092
3 7 609 0 0 4224 0 510 535 0 0 2
649 1080
551 1080
2 6 610 0 0 4224 0 510 535 0 0 2
649 1068
551 1068
1 5 611 0 0 4224 0 510 535 0 0 2
649 1056
551 1056
42
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 40
14 957 187 1021
24 965 176 1013
40 Ligue o "Auto" para 
iniciar a contagem
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 526
1246 162 1659 666
1256 170 1648 570
526 TEMPORIZADOR de 4 bits
0000 
0001
0010
0011 - Usa os 4 primeiros bits de tempo para 
liberar informa��o

0100 
0101 - Ler e decodificar a informa��o

Se for informa��o especial os proximos bits do 
temporizador v�o realizar as sequencias a seguir, 
caso contrario n�o faz nada.

0110
0111 - Pega a e libera a informa��o da proxima 
palavrae coloca em um flip-flop.

1000
1001
1010 - Inseri a infoma��o no lugar que a fun��o 
especial solicitou

1011 - Incrementa o contador e zera o 
temporizador
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 319
-20 1802 261 2207
30 1842 210 2142
319 Tabela de OPCODE

OPCODE - MNEM�NICO 

0000 - MOV A, B
0001 - MOV B, C
0010 - MOV C, A
0011 - ADD A, B
0100 - ADD B, C
0101 - ADD C, A
0110 - AND A, B
0111 - AND B, C
1000 - AND C, A
1001 - OR A, B
1010 - OR B, C
1011 - XOR A, B
1100 - XOR B, C
1101 - LOAD(LD) A
1110 - STORE(ST) A
1111 - DESVIO(JMP)
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
1433 2001 1462 2025
1443 2009 1451 2025
1 B
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
1767 1999 1796 2023
1777 2007 1785 2023
1 C
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 18
1222 951 1387 975
1232 959 1376 975
18 SELETOR DA MEMORIA
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
936 1012 981 1036
946 1020 970 1036
3 REM
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
546 1397 583 1421
556 1405 572 1421
2 RI
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
501 1010 538 1034
511 1018 527 1034
2 PC
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 16
2702 400 2851 424
2712 408 2840 424
16 Menor Relevancia
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 9
1927 740 2020 764
1937 748 2009 764
9 Palavra 1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 9
2210 742 2303 766
2220 750 2292 766
9 Palavra 2
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 9
2503 742 2596 766
2513 750 2585 766
9 Palavra 3
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 9
2808 740 2901 764
2818 748 2890 764
9 Palavra 4
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 9
1926 962 2019 986
1936 970 2008 986
9 Palavra 5
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 9
2211 961 2304 985
2221 969 2293 985
9 Palavra 6
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 9
2503 962 2596 986
2513 970 2585 986
9 Palavra 7
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 9
2806 962 2899 986
2816 970 2888 986
9 Palavra 8
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 9
1926 1176 2019 1200
1936 1184 2008 1200
9 Palavra 9
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 9
2213 1178 2306 1202
2223 1186 2295 1202
9 Palavra10
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 9
2505 1179 2598 1203
2515 1187 2587 1203
9 Palavra11
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 9
2807 1179 2900 1203
2817 1187 2889 1203
9 Palavra12
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 9
1928 1411 2021 1435
1938 1419 2010 1435
9 Palavra13
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 9
2210 1413 2303 1437
2220 1421 2292 1437
9 Palavra14
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 9
2506 1412 2599 1436
2516 1420 2588 1436
9 Palavra15
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 9
2808 1412 2901 1436
2818 1420 2890 1436
9 Palavra16
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
3096 1694 3141 1718
3106 1702 3130 1718
3 RDM
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 79
678 1112 955 1176
688 1120 944 1168
79 Para inserir valores manualmente
basta ligar o logic switch 
"Manual" para 1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 22
731 1088 928 1112
741 1096 917 1112
22 BARRAMENTO DE ENDERE�O
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
1085 1995 1114 2019
1095 2003 1103 2019
1 A
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
2015 1826 2044 1850
2025 1834 2033 1850
1 A
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
2016 1988 2045 2012
2026 1996 2034 2012
1 B
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
2014 2128 2043 2152
2024 2136 2032 2152
1 C
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
2247 1805 2292 1829
2257 1813 2281 1829
3 A+B
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
2248 1964 2293 1988
2258 1972 2282 1988
3 B+C
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
2248 2130 2293 2154
2258 2138 2282 2154
3 C+A
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 33
2879 1917 3076 1961
2889 1925 3065 1957
33 RESPOSTA DAS OPERA��ES 
LOGICAS
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 179
27 1683 264 1847
37 1691 253 1819
179 COLOCAR OS VALORES ANTES DE 
REALIZAR AS OPERA��ES !!!

O INPUT "SET1" quando � 
desativado ativa a opera��o
1 o INPUT "OP" desativa 
todas as opera��es quando
tem valor 1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 106
763 1625 936 1789
773 1633 925 1761
106 Tabela para inserir 
valores manualmente 
para A, B e C

00 pra A
01 pra B
10 pra C
11 n�o faz nada
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 53
78 273 459 317
88 281 448 313
53 CONTADOR DE 0 a 15 Com op��o de incrementar 1 
ou 2
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 16
1770 391 1919 415
1780 399 1908 415
16 Maior Relevancia
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 11
1066 1013 1175 1037
1076 1021 1164 1037
11 Reduz pra 1
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
